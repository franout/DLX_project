
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity complement2_N17_DW01_inc_0 is

   port( A : in std_logic_vector (16 downto 0);  SUM : out std_logic_vector (16
         downto 0));

end complement2_N17_DW01_inc_0;

architecture SYN_rpl of complement2_N17_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port : std_logic;

begin
   
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_16_port, B => A(16), Z => SUM(16));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_1;

architecture SYN_rpl of fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_30_port, SUM_29_port, SUM_28_port, 
      SUM_27_port, SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, 
      SUM_22_port, SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, 
      SUM_17_port, SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, 
      SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port
      , SUM_6_port, SUM_5_port, SUM_4_port, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U2 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U3 : XOR2_X1 port map( A => A(30), B => n56, Z => SUM_30_port);
   U4 : XOR2_X1 port map( A => A(29), B => n55, Z => SUM_29_port);
   U5 : XOR2_X1 port map( A => A(28), B => n54, Z => SUM_28_port);
   U6 : XOR2_X1 port map( A => A(27), B => n53, Z => SUM_27_port);
   U7 : XOR2_X1 port map( A => A(26), B => n52, Z => SUM_26_port);
   U8 : XOR2_X1 port map( A => A(25), B => n51, Z => SUM_25_port);
   U9 : XOR2_X1 port map( A => A(24), B => n50, Z => SUM_24_port);
   U10 : XOR2_X1 port map( A => A(23), B => n49, Z => SUM_23_port);
   U11 : XOR2_X1 port map( A => A(22), B => n48, Z => SUM_22_port);
   U12 : XOR2_X1 port map( A => A(21), B => n47, Z => SUM_21_port);
   U13 : XOR2_X1 port map( A => A(20), B => n46, Z => SUM_20_port);
   U14 : XOR2_X1 port map( A => A(19), B => n45, Z => SUM_19_port);
   U15 : XOR2_X1 port map( A => A(18), B => n44, Z => SUM_18_port);
   U16 : XOR2_X1 port map( A => A(17), B => n43, Z => SUM_17_port);
   U17 : XOR2_X1 port map( A => A(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => A(15), B => n41, Z => SUM_15_port);
   U19 : XOR2_X1 port map( A => A(14), B => n40, Z => SUM_14_port);
   U20 : XOR2_X1 port map( A => A(13), B => n39, Z => SUM_13_port);
   U21 : XOR2_X1 port map( A => A(12), B => n38, Z => SUM_12_port);
   U22 : XOR2_X1 port map( A => A(11), B => n37, Z => SUM_11_port);
   U23 : XOR2_X1 port map( A => A(10), B => n36, Z => SUM_10_port);
   U24 : XOR2_X1 port map( A => A(9), B => n35, Z => SUM_9_port);
   U25 : XOR2_X1 port map( A => A(8), B => n34, Z => SUM_8_port);
   U26 : XOR2_X1 port map( A => A(7), B => n33, Z => SUM_7_port);
   U27 : XOR2_X1 port map( A => A(6), B => n32, Z => SUM_6_port);
   U28 : XOR2_X1 port map( A => A(5), B => n31, Z => SUM_5_port);
   U29 : XOR2_X1 port map( A => A(4), B => n30, Z => SUM_4_port);
   U30 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U31 : NAND2_X1 port map( A1 => A(30), A2 => n56, ZN => n57);
   U32 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n30);
   U33 : AND2_X1 port map( A1 => A(4), A2 => n30, ZN => n31);
   U34 : AND2_X1 port map( A1 => A(5), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => A(6), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => A(7), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => A(8), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => A(9), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => A(10), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => A(11), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => A(12), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => A(13), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => A(14), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => A(15), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => A(16), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => A(17), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => A(18), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => A(19), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => A(20), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => A(21), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => A(22), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => A(23), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => A(24), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => A(25), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => A(26), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => A(27), A2 => n53, ZN => n54);
   U57 : AND2_X1 port map( A1 => A(28), A2 => n54, ZN => n55);
   U58 : AND2_X1 port map( A1 => A(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_0;

architecture SYN_rpl of fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_2_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, SUM_31_port, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => B(2), B => A(2), Z => SUM_2_port);
   U2 : XOR2_X1 port map( A => A(3), B => n31, Z => SUM_3_port);
   U3 : XOR2_X1 port map( A => A(4), B => n32, Z => SUM_4_port);
   U4 : XOR2_X1 port map( A => A(5), B => n33, Z => SUM_5_port);
   U5 : XOR2_X1 port map( A => A(6), B => n34, Z => SUM_6_port);
   U6 : XOR2_X1 port map( A => A(7), B => n35, Z => SUM_7_port);
   U7 : XOR2_X1 port map( A => A(8), B => n36, Z => SUM_8_port);
   U8 : XOR2_X1 port map( A => A(9), B => n37, Z => SUM_9_port);
   U9 : XOR2_X1 port map( A => A(10), B => n38, Z => SUM_10_port);
   U10 : XOR2_X1 port map( A => A(11), B => n39, Z => SUM_11_port);
   U11 : XOR2_X1 port map( A => A(12), B => n40, Z => SUM_12_port);
   U12 : XOR2_X1 port map( A => A(13), B => n41, Z => SUM_13_port);
   U13 : XOR2_X1 port map( A => A(14), B => n42, Z => SUM_14_port);
   U14 : XOR2_X1 port map( A => A(15), B => n43, Z => SUM_15_port);
   U15 : XOR2_X1 port map( A => A(16), B => n44, Z => SUM_16_port);
   U16 : XOR2_X1 port map( A => A(17), B => n45, Z => SUM_17_port);
   U17 : XOR2_X1 port map( A => A(18), B => n46, Z => SUM_18_port);
   U18 : XOR2_X1 port map( A => A(19), B => n47, Z => SUM_19_port);
   U19 : XOR2_X1 port map( A => A(20), B => n48, Z => SUM_20_port);
   U20 : XOR2_X1 port map( A => A(21), B => n49, Z => SUM_21_port);
   U21 : XOR2_X1 port map( A => A(22), B => n50, Z => SUM_22_port);
   U22 : XOR2_X1 port map( A => A(23), B => n51, Z => SUM_23_port);
   U23 : XOR2_X1 port map( A => A(24), B => n52, Z => SUM_24_port);
   U24 : XOR2_X1 port map( A => A(25), B => n53, Z => SUM_25_port);
   U25 : XOR2_X1 port map( A => A(26), B => n54, Z => SUM_26_port);
   U26 : XOR2_X1 port map( A => A(27), B => n55, Z => SUM_27_port);
   U27 : XOR2_X1 port map( A => A(28), B => n56, Z => SUM_28_port);
   U28 : XOR2_X1 port map( A => A(29), B => n57, Z => SUM_29_port);
   U29 : XOR2_X1 port map( A => A(30), B => n58, Z => SUM_30_port);
   U30 : XOR2_X1 port map( A => A(31), B => n59, Z => SUM_31_port);
   U31 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n31);
   U32 : AND2_X1 port map( A1 => A(3), A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => A(4), A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => A(5), A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => A(6), A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => A(7), A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => A(8), A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => A(9), A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => A(10), A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => A(11), A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => A(12), A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => A(13), A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => A(14), A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => A(15), A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => A(16), A2 => n44, ZN => n45);
   U46 : AND2_X1 port map( A1 => A(17), A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => A(18), A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => A(19), A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => A(20), A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => A(21), A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => A(22), A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => A(23), A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => A(24), A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => A(25), A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => A(26), A2 => n54, ZN => n55);
   U56 : AND2_X1 port map( A1 => A(27), A2 => n55, ZN => n56);
   U57 : AND2_X1 port map( A1 => A(28), A2 => n56, ZN => n57);
   U58 : AND2_X1 port map( A1 => A(29), A2 => n57, ZN => n58);
   U59 : AND2_X1 port map( A1 => A(30), A2 => n58, ZN => n59);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT19_DW01_add_0 is

   port( A, B : in std_logic_vector (19 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (19 downto 0);  CO : out std_logic);

end adder_NBIT19_DW01_add_0;

architecture SYN_rpl of adder_NBIT19_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_19_port, carry_18_port, carry_17_port, carry_16_port, 
      carry_15_port, carry_14_port, carry_13_port, carry_12_port, carry_11_port
      , carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      n_1068 : std_logic;

begin
   
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           n_1068, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT21_DW01_add_0 is

   port( A, B : in std_logic_vector (21 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (21 downto 0);  CO : out std_logic);

end adder_NBIT21_DW01_add_0;

architecture SYN_rpl of adder_NBIT21_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_21_port, carry_20_port, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_15_port, carry_14_port, carry_13_port
      , carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port
      , carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, n_1070 : std_logic;

begin
   
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           n_1070, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT23_DW01_add_0 is

   port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (23 downto 0);  CO : out std_logic);

end adder_NBIT23_DW01_add_0;

architecture SYN_rpl of adder_NBIT23_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_23_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, carry_17_port, carry_16_port, carry_15_port
      , carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      n_1072 : std_logic;

begin
   
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           n_1072, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT25_DW01_add_0 is

   port( A, B : in std_logic_vector (25 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (25 downto 0);  CO : out std_logic);

end adder_NBIT25_DW01_add_0;

architecture SYN_rpl of adder_NBIT25_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, n_1074 : std_logic;

begin
   
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           n_1074, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT27_DW01_add_0 is

   port( A, B : in std_logic_vector (27 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (27 downto 0);  CO : out std_logic);

end adder_NBIT27_DW01_add_0;

architecture SYN_rpl of adder_NBIT27_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1076 : 
      std_logic;

begin
   
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           n_1076, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT29_DW01_add_0 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end adder_NBIT29_DW01_add_0;

architecture SYN_rpl of adder_NBIT29_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_29_port, carry_28_port, carry_27_port, carry_26_port, 
      carry_25_port, carry_24_port, carry_23_port, carry_22_port, carry_21_port
      , carry_20_port, carry_19_port, carry_18_port, carry_17_port, 
      carry_16_port, carry_15_port, carry_14_port, carry_13_port, carry_12_port
      , carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port,
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, n_1078 : std_logic;

begin
   
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           n_1078, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT31_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end adder_NBIT31_DW01_add_0;

architecture SYN_rpl of adder_NBIT31_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1080 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1080, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32_DW01_cmp6_1 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end general_alu_N32_DW01_cmp6_1;

architecture SYN_rpl of general_alu_N32_DW01_cmp6_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n69, ZN => n3);
   U2 : INV_X1 port map( A => n129, ZN => n33);
   U3 : INV_X1 port map( A => n117, ZN => n27);
   U4 : INV_X1 port map( A => n93, ZN => n15);
   U5 : INV_X1 port map( A => n81, ZN => n9);
   U6 : INV_X1 port map( A => n105, ZN => n21);
   U7 : INV_X1 port map( A => n132, ZN => n34);
   U8 : INV_X1 port map( A => n120, ZN => n28);
   U9 : INV_X1 port map( A => n108, ZN => n22);
   U10 : INV_X1 port map( A => n96, ZN => n16);
   U11 : INV_X1 port map( A => n84, ZN => n10);
   U12 : INV_X1 port map( A => n72, ZN => n4);
   U13 : INV_X1 port map( A => n144, ZN => n40);
   U14 : INV_X1 port map( A => n142, ZN => n36);
   U15 : INV_X1 port map( A => n145, ZN => n38);
   U16 : INV_X1 port map( A => n118, ZN => n24);
   U17 : INV_X1 port map( A => n121, ZN => n26);
   U18 : INV_X1 port map( A => n94, ZN => n12);
   U19 : INV_X1 port map( A => n97, ZN => n14);
   U20 : INV_X1 port map( A => n130, ZN => n30);
   U21 : INV_X1 port map( A => n82, ZN => n6);
   U22 : INV_X1 port map( A => n106, ZN => n18);
   U23 : INV_X1 port map( A => n70, ZN => n1);
   U24 : INV_X1 port map( A => n73, ZN => n2);
   U25 : INV_X1 port map( A => n133, ZN => n32);
   U26 : INV_X1 port map( A => n85, ZN => n8);
   U27 : INV_X1 port map( A => n109, ZN => n20);
   U28 : INV_X1 port map( A => n141, ZN => n39);
   U29 : INV_X1 port map( A => n152, ZN => n44);
   U30 : INV_X1 port map( A => n201, ZN => n43);
   U31 : INV_X1 port map( A => B(4), ZN => n41);
   U32 : INV_X1 port map( A => B(8), ZN => n35);
   U33 : INV_X1 port map( A => B(16), ZN => n23);
   U34 : INV_X1 port map( A => B(20), ZN => n17);
   U35 : INV_X1 port map( A => B(24), ZN => n11);
   U36 : INV_X1 port map( A => B(14), ZN => n25);
   U37 : INV_X1 port map( A => B(6), ZN => n37);
   U38 : INV_X1 port map( A => B(10), ZN => n31);
   U39 : INV_X1 port map( A => B(12), ZN => n29);
   U40 : INV_X1 port map( A => B(18), ZN => n19);
   U41 : INV_X1 port map( A => B(22), ZN => n13);
   U42 : INV_X1 port map( A => B(26), ZN => n7);
   U43 : INV_X1 port map( A => A(1), ZN => n61);
   U44 : INV_X1 port map( A => B(28), ZN => n5);
   U45 : INV_X1 port map( A => B(2), ZN => n42);
   U46 : INV_X1 port map( A => A(0), ZN => n62);
   U47 : INV_X1 port map( A => A(3), ZN => n60);
   U48 : INV_X1 port map( A => A(5), ZN => n59);
   U49 : INV_X1 port map( A => A(13), ZN => n55);
   U50 : INV_X1 port map( A => A(21), ZN => n51);
   U51 : INV_X1 port map( A => A(25), ZN => n49);
   U52 : INV_X1 port map( A => A(9), ZN => n57);
   U53 : INV_X1 port map( A => A(15), ZN => n54);
   U54 : INV_X1 port map( A => A(31), ZN => n45);
   U55 : INV_X1 port map( A => A(17), ZN => n53);
   U56 : INV_X1 port map( A => A(29), ZN => n47);
   U57 : INV_X1 port map( A => A(11), ZN => n56);
   U58 : INV_X1 port map( A => A(27), ZN => n48);
   U59 : INV_X1 port map( A => A(19), ZN => n52);
   U60 : INV_X1 port map( A => A(23), ZN => n50);
   U61 : INV_X1 port map( A => A(7), ZN => n58);
   U62 : INV_X1 port map( A => A(30), ZN => n46);
   U63 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => LE);
   U64 : NAND3_X1 port map( A1 => n65, A2 => n66, A3 => n67, ZN => n64);
   U65 : NAND3_X1 port map( A1 => n68, A2 => n69, A3 => n1, ZN => n65);
   U66 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n2, ZN => n68);
   U67 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => n71);
   U68 : NAND3_X1 port map( A1 => n77, A2 => n78, A3 => n79, ZN => n74);
   U69 : NAND3_X1 port map( A1 => n80, A2 => n81, A3 => n6, ZN => n77);
   U70 : NAND3_X1 port map( A1 => n83, A2 => n84, A3 => n8, ZN => n80);
   U71 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => n83);
   U72 : NAND3_X1 port map( A1 => n89, A2 => n90, A3 => n91, ZN => n86);
   U73 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n12, ZN => n89);
   U74 : NAND3_X1 port map( A1 => n95, A2 => n96, A3 => n14, ZN => n92);
   U75 : NAND3_X1 port map( A1 => n98, A2 => n99, A3 => n100, ZN => n95);
   U76 : NAND3_X1 port map( A1 => n101, A2 => n102, A3 => n103, ZN => n98);
   U77 : NAND3_X1 port map( A1 => n104, A2 => n105, A3 => n18, ZN => n101);
   U78 : NAND3_X1 port map( A1 => n107, A2 => n108, A3 => n20, ZN => n104);
   U79 : NAND3_X1 port map( A1 => n110, A2 => n111, A3 => n112, ZN => n107);
   U80 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n115, ZN => n110);
   U81 : NAND3_X1 port map( A1 => n116, A2 => n117, A3 => n24, ZN => n113);
   U82 : NAND3_X1 port map( A1 => n119, A2 => n120, A3 => n26, ZN => n116);
   U83 : NAND3_X1 port map( A1 => n122, A2 => n123, A3 => n124, ZN => n119);
   U84 : NAND3_X1 port map( A1 => n125, A2 => n126, A3 => n127, ZN => n122);
   U85 : NAND3_X1 port map( A1 => n128, A2 => n129, A3 => n30, ZN => n125);
   U86 : NAND3_X1 port map( A1 => n131, A2 => n132, A3 => n32, ZN => n128);
   U87 : NAND3_X1 port map( A1 => n134, A2 => n135, A3 => n136, ZN => n131);
   U88 : NAND3_X1 port map( A1 => n137, A2 => n138, A3 => n139, ZN => n134);
   U89 : NAND3_X1 port map( A1 => n140, A2 => n141, A3 => n36, ZN => n137);
   U90 : NAND3_X1 port map( A1 => n143, A2 => n144, A3 => n38, ZN => n140);
   U91 : NAND3_X1 port map( A1 => n146, A2 => n147, A3 => n148, ZN => n143);
   U92 : NAND3_X1 port map( A1 => n149, A2 => n150, A3 => n151, ZN => n146);
   U93 : OAI211_X1 port map( C1 => A(1), C2 => n152, A => n153, B => n154, ZN 
                           => n149);
   U94 : OAI21_X1 port map( B1 => n44, B2 => n61, A => B(1), ZN => n153);
   U95 : NOR2_X1 port map( A1 => n62, A2 => B(0), ZN => n152);
   U96 : OAI21_X1 port map( B1 => n155, B2 => n156, A => n67, ZN => GE);
   U97 : NAND2_X1 port map( A1 => B(31), A2 => n45, ZN => n67);
   U98 : NAND2_X1 port map( A1 => n63, A2 => n157, ZN => n156);
   U99 : OR2_X1 port map( A1 => n45, A2 => B(31), ZN => n63);
   U100 : AOI211_X1 port map( C1 => n158, C2 => n159, A => n70, B => n73, ZN =>
                           n155);
   U101 : NOR2_X1 port map( A1 => n47, A2 => B(29), ZN => n73);
   U102 : NAND2_X1 port map( A1 => n66, A2 => n157, ZN => n70);
   U103 : NAND2_X1 port map( A1 => B(30), A2 => n46, ZN => n157);
   U104 : OR2_X1 port map( A1 => n46, A2 => B(30), ZN => n66);
   U105 : OAI211_X1 port map( C1 => n160, C2 => n161, A => n79, B => n76, ZN =>
                           n159);
   U106 : NOR2_X1 port map( A1 => n162, A2 => n4, ZN => n76);
   U107 : NAND2_X1 port map( A1 => A(28), A2 => n5, ZN => n72);
   U108 : OR2_X1 port map( A1 => n48, A2 => B(27), ZN => n79);
   U109 : NAND2_X1 port map( A1 => n75, A2 => n163, ZN => n161);
   U110 : NAND2_X1 port map( A1 => B(27), A2 => n48, ZN => n75);
   U111 : AOI211_X1 port map( C1 => n164, C2 => n165, A => n82, B => n85, ZN =>
                           n160);
   U112 : NOR2_X1 port map( A1 => n49, A2 => B(25), ZN => n85);
   U113 : NAND2_X1 port map( A1 => n163, A2 => n78, ZN => n82);
   U114 : NAND2_X1 port map( A1 => A(26), A2 => n7, ZN => n78);
   U115 : OR2_X1 port map( A1 => n7, A2 => A(26), ZN => n163);
   U116 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n91, B => n88, ZN =>
                           n165);
   U117 : NOR2_X1 port map( A1 => n168, A2 => n10, ZN => n88);
   U118 : NAND2_X1 port map( A1 => A(24), A2 => n11, ZN => n84);
   U119 : OR2_X1 port map( A1 => n50, A2 => B(23), ZN => n91);
   U120 : NAND2_X1 port map( A1 => n87, A2 => n169, ZN => n167);
   U121 : NAND2_X1 port map( A1 => B(23), A2 => n50, ZN => n87);
   U122 : AOI211_X1 port map( C1 => n170, C2 => n171, A => n94, B => n97, ZN =>
                           n166);
   U123 : NOR2_X1 port map( A1 => n51, A2 => B(21), ZN => n97);
   U124 : NAND2_X1 port map( A1 => n169, A2 => n90, ZN => n94);
   U125 : NAND2_X1 port map( A1 => A(22), A2 => n13, ZN => n90);
   U126 : OR2_X1 port map( A1 => n13, A2 => A(22), ZN => n169);
   U127 : OAI211_X1 port map( C1 => n172, C2 => n173, A => n103, B => n100, ZN 
                           => n171);
   U128 : NOR2_X1 port map( A1 => n174, A2 => n16, ZN => n100);
   U129 : NAND2_X1 port map( A1 => A(20), A2 => n17, ZN => n96);
   U130 : OR2_X1 port map( A1 => n52, A2 => B(19), ZN => n103);
   U131 : NAND2_X1 port map( A1 => n99, A2 => n175, ZN => n173);
   U132 : NAND2_X1 port map( A1 => B(19), A2 => n52, ZN => n99);
   U133 : AOI211_X1 port map( C1 => n176, C2 => n177, A => n106, B => n109, ZN 
                           => n172);
   U134 : NOR2_X1 port map( A1 => n53, A2 => B(17), ZN => n109);
   U135 : NAND2_X1 port map( A1 => n175, A2 => n102, ZN => n106);
   U136 : NAND2_X1 port map( A1 => A(18), A2 => n19, ZN => n102);
   U137 : OR2_X1 port map( A1 => n19, A2 => A(18), ZN => n175);
   U138 : OAI211_X1 port map( C1 => n178, C2 => n179, A => n115, B => n112, ZN 
                           => n177);
   U139 : NOR2_X1 port map( A1 => n180, A2 => n22, ZN => n112);
   U140 : NAND2_X1 port map( A1 => A(16), A2 => n23, ZN => n108);
   U141 : OR2_X1 port map( A1 => n54, A2 => B(15), ZN => n115);
   U142 : NAND2_X1 port map( A1 => n111, A2 => n181, ZN => n179);
   U143 : NAND2_X1 port map( A1 => B(15), A2 => n54, ZN => n111);
   U144 : AOI211_X1 port map( C1 => n182, C2 => n183, A => n118, B => n121, ZN 
                           => n178);
   U145 : NOR2_X1 port map( A1 => n55, A2 => B(13), ZN => n121);
   U146 : NAND2_X1 port map( A1 => n181, A2 => n114, ZN => n118);
   U147 : NAND2_X1 port map( A1 => A(14), A2 => n25, ZN => n114);
   U148 : OR2_X1 port map( A1 => n25, A2 => A(14), ZN => n181);
   U149 : OAI211_X1 port map( C1 => n184, C2 => n185, A => n127, B => n124, ZN 
                           => n183);
   U150 : NOR2_X1 port map( A1 => n186, A2 => n28, ZN => n124);
   U151 : NAND2_X1 port map( A1 => A(12), A2 => n29, ZN => n120);
   U152 : OR2_X1 port map( A1 => n56, A2 => B(11), ZN => n127);
   U153 : NAND2_X1 port map( A1 => n123, A2 => n187, ZN => n185);
   U154 : NAND2_X1 port map( A1 => B(11), A2 => n56, ZN => n123);
   U155 : AOI211_X1 port map( C1 => n188, C2 => n189, A => n130, B => n133, ZN 
                           => n184);
   U156 : NOR2_X1 port map( A1 => n57, A2 => B(9), ZN => n133);
   U157 : NAND2_X1 port map( A1 => n187, A2 => n126, ZN => n130);
   U158 : NAND2_X1 port map( A1 => A(10), A2 => n31, ZN => n126);
   U159 : OR2_X1 port map( A1 => n31, A2 => A(10), ZN => n187);
   U160 : OAI211_X1 port map( C1 => n190, C2 => n191, A => n139, B => n136, ZN 
                           => n189);
   U161 : NOR2_X1 port map( A1 => n192, A2 => n34, ZN => n136);
   U162 : NAND2_X1 port map( A1 => A(8), A2 => n35, ZN => n132);
   U163 : OR2_X1 port map( A1 => n58, A2 => B(7), ZN => n139);
   U164 : NAND2_X1 port map( A1 => n135, A2 => n193, ZN => n191);
   U165 : NAND2_X1 port map( A1 => B(7), A2 => n58, ZN => n135);
   U166 : AOI211_X1 port map( C1 => n194, C2 => n195, A => n142, B => n145, ZN 
                           => n190);
   U167 : NOR2_X1 port map( A1 => n59, A2 => B(5), ZN => n145);
   U168 : NAND2_X1 port map( A1 => n193, A2 => n138, ZN => n142);
   U169 : NAND2_X1 port map( A1 => A(6), A2 => n37, ZN => n138);
   U170 : OR2_X1 port map( A1 => n37, A2 => A(6), ZN => n193);
   U171 : NAND3_X1 port map( A1 => n196, A2 => n151, A3 => n148, ZN => n195);
   U172 : NOR2_X1 port map( A1 => n197, A2 => n40, ZN => n148);
   U173 : NAND2_X1 port map( A1 => A(4), A2 => n41, ZN => n144);
   U174 : OR2_X1 port map( A1 => n60, A2 => B(3), ZN => n151);
   U175 : NAND3_X1 port map( A1 => n147, A2 => n198, A3 => n199, ZN => n196);
   U176 : OAI211_X1 port map( C1 => n200, C2 => n61, A => n43, B => n154, ZN =>
                           n199);
   U177 : AND2_X1 port map( A1 => n198, A2 => n150, ZN => n154);
   U178 : NAND2_X1 port map( A1 => A(2), A2 => n42, ZN => n150);
   U179 : AOI21_X1 port map( B1 => n61, B2 => n200, A => B(1), ZN => n201);
   U180 : AND2_X1 port map( A1 => B(0), A2 => n62, ZN => n200);
   U181 : OR2_X1 port map( A1 => n42, A2 => A(2), ZN => n198);
   U182 : NAND2_X1 port map( A1 => B(3), A2 => n60, ZN => n147);
   U183 : NOR2_X1 port map( A1 => n197, A2 => n39, ZN => n194);
   U184 : NAND2_X1 port map( A1 => B(5), A2 => n59, ZN => n141);
   U185 : NOR2_X1 port map( A1 => n41, A2 => A(4), ZN => n197);
   U186 : NOR2_X1 port map( A1 => n192, A2 => n33, ZN => n188);
   U187 : NAND2_X1 port map( A1 => B(9), A2 => n57, ZN => n129);
   U188 : NOR2_X1 port map( A1 => n35, A2 => A(8), ZN => n192);
   U189 : NOR2_X1 port map( A1 => n186, A2 => n27, ZN => n182);
   U190 : NAND2_X1 port map( A1 => B(13), A2 => n55, ZN => n117);
   U191 : NOR2_X1 port map( A1 => n29, A2 => A(12), ZN => n186);
   U192 : NOR2_X1 port map( A1 => n180, A2 => n21, ZN => n176);
   U193 : NAND2_X1 port map( A1 => B(17), A2 => n53, ZN => n105);
   U194 : NOR2_X1 port map( A1 => n23, A2 => A(16), ZN => n180);
   U195 : NOR2_X1 port map( A1 => n174, A2 => n15, ZN => n170);
   U196 : NAND2_X1 port map( A1 => B(21), A2 => n51, ZN => n93);
   U197 : NOR2_X1 port map( A1 => n17, A2 => A(20), ZN => n174);
   U198 : NOR2_X1 port map( A1 => n168, A2 => n9, ZN => n164);
   U199 : NAND2_X1 port map( A1 => B(25), A2 => n49, ZN => n81);
   U200 : NOR2_X1 port map( A1 => n11, A2 => A(24), ZN => n168);
   U201 : NOR2_X1 port map( A1 => n162, A2 => n3, ZN => n158);
   U202 : NAND2_X1 port map( A1 => B(29), A2 => n47, ZN => n69);
   U203 : NOR2_X1 port map( A1 => n5, A2 => A(28), ZN => n162);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end general_alu_N32_DW01_cmp6_0;

architecture SYN_rpl of general_alu_N32_DW01_cmp6_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B(1), ZN => n2);
   U2 : INV_X1 port map( A => A(1), ZN => n1);
   U3 : INV_X1 port map( A => B(0), ZN => n3);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => NE);
   U5 : NOR4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U6 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => n9
                           );
   U7 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n13);
   U8 : XNOR2_X1 port map( A => B(13), B => A(13), ZN => n12);
   U9 : XNOR2_X1 port map( A => B(14), B => A(14), ZN => n11);
   U10 : XNOR2_X1 port map( A => B(15), B => A(15), ZN => n10);
   U11 : NAND4_X1 port map( A1 => n14, A2 => n15, A3 => n16, A4 => n17, ZN => 
                           n8);
   U12 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n17);
   U13 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n16);
   U14 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n15);
   U15 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n14);
   U16 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n7);
   U17 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n21);
   U18 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n20);
   U19 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n19);
   U20 : XNOR2_X1 port map( A => B(7), B => A(7), ZN => n18);
   U21 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           n6);
   U22 : OAI22_X1 port map( A1 => A(1), A2 => n26, B1 => n26, B2 => n2, ZN => 
                           n25);
   U23 : AND2_X1 port map( A1 => A(0), A2 => n3, ZN => n26);
   U24 : OAI22_X1 port map( A1 => n27, A2 => n1, B1 => B(1), B2 => n27, ZN => 
                           n24);
   U25 : NOR2_X1 port map( A1 => n3, A2 => A(0), ZN => n27);
   U26 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n23);
   U27 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n22);
   U28 : NOR4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => n4
                           );
   U29 : NAND4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => 
                           n31);
   U30 : XNOR2_X1 port map( A => B(28), B => A(28), ZN => n35);
   U31 : XNOR2_X1 port map( A => B(29), B => A(29), ZN => n34);
   U32 : XNOR2_X1 port map( A => B(30), B => A(30), ZN => n33);
   U33 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n32);
   U34 : NAND4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => 
                           n30);
   U35 : XNOR2_X1 port map( A => B(24), B => A(24), ZN => n39);
   U36 : XNOR2_X1 port map( A => B(25), B => A(25), ZN => n38);
   U37 : XNOR2_X1 port map( A => B(26), B => A(26), ZN => n37);
   U38 : XNOR2_X1 port map( A => B(27), B => A(27), ZN => n36);
   U39 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n29);
   U40 : XNOR2_X1 port map( A => B(20), B => A(20), ZN => n43);
   U41 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n42);
   U42 : XNOR2_X1 port map( A => B(22), B => A(22), ZN => n41);
   U43 : XNOR2_X1 port map( A => B(23), B => A(23), ZN => n40);
   U44 : NAND4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => 
                           n28);
   U45 : XNOR2_X1 port map( A => B(16), B => A(16), ZN => n47);
   U46 : XNOR2_X1 port map( A => B(17), B => A(17), ZN => n46);
   U47 : XNOR2_X1 port map( A => B(18), B => A(18), ZN => n45);
   U48 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => n44);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_7 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_7;

architecture SYN_STRUCTURAL of RCA_NBIT8_7 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_52 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_51 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_50 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_49 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_6 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_6;

architecture SYN_STRUCTURAL of RCA_NBIT8_6 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_44 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_43 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_42 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_41 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_5 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_5;

architecture SYN_STRUCTURAL of RCA_NBIT8_5 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_36 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_35 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_34 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_33 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_4 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_4;

architecture SYN_STRUCTURAL of RCA_NBIT8_4 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_28 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_27 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_26 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_25 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_3 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_3;

architecture SYN_STRUCTURAL of RCA_NBIT8_3 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_20 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_19 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_18 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_17 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_2 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_2;

architecture SYN_STRUCTURAL of RCA_NBIT8_2 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_12 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_11 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_10 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_9 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_1 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_1;

architecture SYN_STRUCTURAL of RCA_NBIT8_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_4 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_3 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_2 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_1 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT8_3 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0));

end CSB_NBIT8_3;

architecture SYN_STRUCTURAL of CSB_NBIT8_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_NBIT8_5
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT8_6
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_c0_7_port, out_c0_6_port, 
      out_c0_5_port, out_c0_4_port, out_c0_3_port, out_c0_2_port, out_c0_1_port
      , out_c0_0_port, out_c1_7_port, out_c1_6_port, out_c1_5_port, 
      out_c1_4_port, out_c1_3_port, out_c1_2_port, out_c1_1_port, out_c1_0_port
      , n_1092, n_1093 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT8_6 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(7) => 
                           out_c0_7_port, S(6) => out_c0_6_port, S(5) => 
                           out_c0_5_port, S(4) => out_c0_4_port, S(3) => 
                           out_c0_3_port, S(2) => out_c0_2_port, S(1) => 
                           out_c0_1_port, S(0) => out_c0_0_port, Co => n_1092);
   RCA1 : RCA_NBIT8_5 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(7) => 
                           out_c1_7_port, S(6) => out_c1_6_port, S(5) => 
                           out_c1_5_port, S(4) => out_c1_4_port, S(3) => 
                           out_c1_3_port, S(2) => out_c1_2_port, S(1) => 
                           out_c1_1_port, S(0) => out_c1_0_port, Co => n_1093);
   U3 : MUX2_X1 port map( A => out_c0_7_port, B => out_c1_7_port, S => Ci, Z =>
                           S(7));
   U4 : MUX2_X1 port map( A => out_c0_6_port, B => out_c1_6_port, S => Ci, Z =>
                           S(6));
   U5 : MUX2_X1 port map( A => out_c0_5_port, B => out_c1_5_port, S => Ci, Z =>
                           S(5));
   U6 : MUX2_X1 port map( A => out_c0_4_port, B => out_c1_4_port, S => Ci, Z =>
                           S(4));
   U7 : MUX2_X1 port map( A => out_c0_3_port, B => out_c1_3_port, S => Ci, Z =>
                           S(3));
   U8 : MUX2_X1 port map( A => out_c0_2_port, B => out_c1_2_port, S => Ci, Z =>
                           S(2));
   U9 : MUX2_X1 port map( A => out_c0_1_port, B => out_c1_1_port, S => Ci, Z =>
                           S(1));
   U10 : MUX2_X1 port map( A => out_c0_0_port, B => out_c1_0_port, S => Ci, Z 
                           => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT8_2 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0));

end CSB_NBIT8_2;

architecture SYN_STRUCTURAL of CSB_NBIT8_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_NBIT8_3
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT8_4
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_c0_7_port, out_c0_6_port, 
      out_c0_5_port, out_c0_4_port, out_c0_3_port, out_c0_2_port, out_c0_1_port
      , out_c0_0_port, out_c1_7_port, out_c1_6_port, out_c1_5_port, 
      out_c1_4_port, out_c1_3_port, out_c1_2_port, out_c1_1_port, out_c1_0_port
      , n_1094, n_1095 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT8_4 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(7) => 
                           out_c0_7_port, S(6) => out_c0_6_port, S(5) => 
                           out_c0_5_port, S(4) => out_c0_4_port, S(3) => 
                           out_c0_3_port, S(2) => out_c0_2_port, S(1) => 
                           out_c0_1_port, S(0) => out_c0_0_port, Co => n_1094);
   RCA1 : RCA_NBIT8_3 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(7) => 
                           out_c1_7_port, S(6) => out_c1_6_port, S(5) => 
                           out_c1_5_port, S(4) => out_c1_4_port, S(3) => 
                           out_c1_3_port, S(2) => out_c1_2_port, S(1) => 
                           out_c1_1_port, S(0) => out_c1_0_port, Co => n_1095);
   U3 : MUX2_X1 port map( A => out_c0_7_port, B => out_c1_7_port, S => Ci, Z =>
                           S(7));
   U4 : MUX2_X1 port map( A => out_c0_6_port, B => out_c1_6_port, S => Ci, Z =>
                           S(6));
   U5 : MUX2_X1 port map( A => out_c0_5_port, B => out_c1_5_port, S => Ci, Z =>
                           S(5));
   U6 : MUX2_X1 port map( A => out_c0_4_port, B => out_c1_4_port, S => Ci, Z =>
                           S(4));
   U7 : MUX2_X1 port map( A => out_c0_3_port, B => out_c1_3_port, S => Ci, Z =>
                           S(3));
   U8 : MUX2_X1 port map( A => out_c0_2_port, B => out_c1_2_port, S => Ci, Z =>
                           S(2));
   U9 : MUX2_X1 port map( A => out_c0_1_port, B => out_c1_1_port, S => Ci, Z =>
                           S(1));
   U10 : MUX2_X1 port map( A => out_c0_0_port, B => out_c1_0_port, S => Ci, Z 
                           => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT8_1 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0));

end CSB_NBIT8_1;

architecture SYN_STRUCTURAL of CSB_NBIT8_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_NBIT8_1
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT8_2
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_c0_7_port, out_c0_6_port, 
      out_c0_5_port, out_c0_4_port, out_c0_3_port, out_c0_2_port, out_c0_1_port
      , out_c0_0_port, out_c1_7_port, out_c1_6_port, out_c1_5_port, 
      out_c1_4_port, out_c1_3_port, out_c1_2_port, out_c1_1_port, out_c1_0_port
      , n_1096, n_1097 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT8_2 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(7) => 
                           out_c0_7_port, S(6) => out_c0_6_port, S(5) => 
                           out_c0_5_port, S(4) => out_c0_4_port, S(3) => 
                           out_c0_3_port, S(2) => out_c0_2_port, S(1) => 
                           out_c0_1_port, S(0) => out_c0_0_port, Co => n_1096);
   RCA1 : RCA_NBIT8_1 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(7) => 
                           out_c1_7_port, S(6) => out_c1_6_port, S(5) => 
                           out_c1_5_port, S(4) => out_c1_4_port, S(3) => 
                           out_c1_3_port, S(2) => out_c1_2_port, S(1) => 
                           out_c1_1_port, S(0) => out_c1_0_port, Co => n_1097);
   U3 : MUX2_X1 port map( A => out_c0_7_port, B => out_c1_7_port, S => Ci, Z =>
                           S(7));
   U4 : MUX2_X1 port map( A => out_c0_6_port, B => out_c1_6_port, S => Ci, Z =>
                           S(6));
   U5 : MUX2_X1 port map( A => out_c0_5_port, B => out_c1_5_port, S => Ci, Z =>
                           S(5));
   U6 : MUX2_X1 port map( A => out_c0_4_port, B => out_c1_4_port, S => Ci, Z =>
                           S(4));
   U7 : MUX2_X1 port map( A => out_c0_3_port, B => out_c1_3_port, S => Ci, Z =>
                           S(3));
   U8 : MUX2_X1 port map( A => out_c0_2_port, B => out_c1_2_port, S => Ci, Z =>
                           S(2));
   U9 : MUX2_X1 port map( A => out_c0_1_port, B => out_c1_1_port, S => Ci, Z =>
                           S(1));
   U10 : MUX2_X1 port map( A => out_c0_0_port, B => out_c1_0_port, S => Ci, Z 
                           => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_26 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_26;

architecture SYN_BEHAVIORAL of PGSB_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_25 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_25;

architecture SYN_BEHAVIORAL of PGSB_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_24 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_24;

architecture SYN_BEHAVIORAL of PGSB_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_23 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_23;

architecture SYN_BEHAVIORAL of PGSB_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_22 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_22;

architecture SYN_BEHAVIORAL of PGSB_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_21 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_21;

architecture SYN_BEHAVIORAL of PGSB_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_20 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_20;

architecture SYN_BEHAVIORAL of PGSB_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_19 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_19;

architecture SYN_BEHAVIORAL of PGSB_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_18 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_18;

architecture SYN_BEHAVIORAL of PGSB_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_17 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_17;

architecture SYN_BEHAVIORAL of PGSB_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_16 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_16;

architecture SYN_BEHAVIORAL of PGSB_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_15 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_15;

architecture SYN_BEHAVIORAL of PGSB_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_14 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_14;

architecture SYN_BEHAVIORAL of PGSB_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_13 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_13;

architecture SYN_BEHAVIORAL of PGSB_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_12 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_12;

architecture SYN_BEHAVIORAL of PGSB_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_11 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_11;

architecture SYN_BEHAVIORAL of PGSB_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_10 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_10;

architecture SYN_BEHAVIORAL of PGSB_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_9 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_9;

architecture SYN_BEHAVIORAL of PGSB_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_8 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_8;

architecture SYN_BEHAVIORAL of PGSB_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_7 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_7;

architecture SYN_BEHAVIORAL of PGSB_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_6 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_6;

architecture SYN_BEHAVIORAL of PGSB_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_5 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_5;

architecture SYN_BEHAVIORAL of PGSB_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_4 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_4;

architecture SYN_BEHAVIORAL of PGSB_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_3 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_3;

architecture SYN_BEHAVIORAL of PGSB_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_2 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_2;

architecture SYN_BEHAVIORAL of PGSB_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_1 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_1;

architecture SYN_BEHAVIORAL of PGSB_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_8 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_8;

architecture SYN_BEHAVIORAL of GSB_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_7 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_7;

architecture SYN_BEHAVIORAL of GSB_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_6 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_6;

architecture SYN_BEHAVIORAL of GSB_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_5 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_5;

architecture SYN_BEHAVIORAL of GSB_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_4 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_4;

architecture SYN_BEHAVIORAL of GSB_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_3 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_3;

architecture SYN_BEHAVIORAL of GSB_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_2 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_2;

architecture SYN_BEHAVIORAL of GSB_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_1 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_1;

architecture SYN_BEHAVIORAL of GSB_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_5 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_5;

architecture SYN_struc of reg_nbit_n16_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_65
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_66
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_67
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_68
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_69
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_70
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_71
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_72
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_73
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_74
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_75
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_76
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_77
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_78
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_79
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_80
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_80 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_79 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_78 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_77 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_76 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_75 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_74 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_73 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_72 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_71 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_70 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_69 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_68 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_67 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_66 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_65 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_4 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_4;

architecture SYN_struc of reg_nbit_n16_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_49
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_50
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_51
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_52
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_53
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_54
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_55
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_56
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_57
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_58
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_59
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_60
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_61
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_62
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_63
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_64
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_64 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_63 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_62 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_61 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_60 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_59 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_58 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_57 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_56 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_55 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_54 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_53 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_52 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_51 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_50 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_49 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_3 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_3;

architecture SYN_struc of reg_nbit_n16_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_33
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_34
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_35
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_36
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_37
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_38
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_39
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_40
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_41
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_42
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_43
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_44
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_45
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_46
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_47
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_48
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_48 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_47 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_46 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_45 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_44 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_43 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_42 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_41 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_40 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_39 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_38 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_37 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_36 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_35 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_34 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_33 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_2 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_2;

architecture SYN_struc of reg_nbit_n16_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_17
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_18
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_19
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_20
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_21
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_22
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_23
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_24
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_25
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_26
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_27
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_28
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_29
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_30
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_31
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_32
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_32 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_31 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_30 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_29 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_28 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_27 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_26 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_25 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_24 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_23 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_22 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_21 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_20 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_19 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_18 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_17 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_1;

architecture SYN_struc of reg_nbit_n16_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_3
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_4
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_5
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_6
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_7
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_8
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_9
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_10
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_11
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_12
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_13
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_14
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_15
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_16
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_16 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_15 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_14 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_13 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_12 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_11 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_10 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_9 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_8 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_7 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_6 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_5 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_4 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_3 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_2 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_1 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_5 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_5;

architecture SYN_struc of reg_nbit_n249_5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1221
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1222
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1223
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1224
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1225
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1226
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1227
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1228
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1229
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1230
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1231
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1232
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1233
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1234
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1235
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1236
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1237
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1238
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1239
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1240
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1241
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1242
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1243
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1244
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1245
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1246
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1247
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1248
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1249
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1250
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1251
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1252
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1253
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1254
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1255
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1256
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1257
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1258
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1259
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1260
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1261
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1262
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1263
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1264
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1265
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1266
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1267
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1268
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1269
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1270
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1271
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1272
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1273
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1274
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1275
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1276
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1277
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1278
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1279
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1280
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1281
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1282
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1283
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1284
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1285
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1286
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1287
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1288
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1289
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1290
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1291
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1292
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1293
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1294
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1295
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1296
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1297
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1298
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1299
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1300
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1301
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1302
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1303
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1304
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1305
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1306
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1307
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1308
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1309
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1310
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1311
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1312
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1313
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1314
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1315
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1316
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1317
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1318
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1319
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1320
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1321
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1322
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1323
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1324
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1325
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1326
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1327
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1328
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1329
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1330
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1331
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1332
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1333
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1334
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1335
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1336
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1337
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1338
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1339
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1340
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1341
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1342
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1343
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1344
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1345
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1346
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1347
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1348
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1349
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1350
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1351
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1352
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1353
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1354
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1355
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1356
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1357
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1358
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1359
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1360
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1361
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1362
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1363
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1364
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1365
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1366
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1367
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1368
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1369
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1370
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1371
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1372
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1373
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1374
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1375
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1376
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1377
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1378
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1379
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1380
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1381
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1382
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1383
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1384
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1385
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1386
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1387
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1388
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1389
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1390
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1391
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1392
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1393
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1394
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1395
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1396
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1397
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1398
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1399
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1400
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1401
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1402
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1403
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1404
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1405
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1406
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1407
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1408
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1409
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1410
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1411
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1412
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1413
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1414
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1415
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1416
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1417
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1418
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1419
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1420
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1421
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1422
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1423
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1424
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1425
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1426
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1427
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1428
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1429
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1430
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1431
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1432
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1433
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1434
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1435
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1436
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1437
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1438
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1439
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1440
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1441
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1442
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1443
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1444
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1445
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1446
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1447
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1448
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1449
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1450
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1451
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1452
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1453
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1454
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1455
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1456
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1457
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1458
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1459
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1460
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1461
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1462
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1463
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1464
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1465
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1466
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1467
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1468
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1469
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_1469 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_1468 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_1467 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_1466 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_1465 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_1464 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_1463 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_1462 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_1461 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_1460 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_1459 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_1458 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_1457 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_1456 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_1455 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_1454 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_1453 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_1452 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_1451 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_1450 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_1449 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_1448 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_1447 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_1446 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_1445 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_1444 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_1443 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_1442 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_1441 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_1440 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_1439 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_1438 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_1437 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_1436 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_1435 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_1434 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_1433 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_1432 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_1431 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_1430 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_1429 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_1428 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_1427 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_1426 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_1425 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_1424 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_1423 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_1422 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_1421 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_1420 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_1419 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_1418 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_1417 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_1416 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_1415 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_1414 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_1413 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_1412 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_1411 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_1410 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_1409 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_1408 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_1407 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_1406 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_1405 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_1404 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_1403 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_1402 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_1401 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_1400 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_1399 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_1398 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_1397 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_1396 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_1395 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_1394 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_1393 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_1392 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_1391 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_1390 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_1389 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_1388 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_1387 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_1386 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_1385 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_1384 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_1383 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_1382 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_1381 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_1380 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_1379 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_1378 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_1377 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_1376 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_1375 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_1374 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_1373 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_1372 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_1371 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_1370 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_1369 port map( D => d(100), CK => n43, RESET => n15, Q => 
                           Q(100));
   D_I_101 : FD_1368 port map( D => d(101), CK => n43, RESET => n15, Q => 
                           Q(101));
   D_I_102 : FD_1367 port map( D => d(102), CK => n43, RESET => n15, Q => 
                           Q(102));
   D_I_103 : FD_1366 port map( D => d(103), CK => n43, RESET => n15, Q => 
                           Q(103));
   D_I_104 : FD_1365 port map( D => d(104), CK => n43, RESET => n15, Q => 
                           Q(104));
   D_I_105 : FD_1364 port map( D => d(105), CK => n43, RESET => n15, Q => 
                           Q(105));
   D_I_106 : FD_1363 port map( D => d(106), CK => n43, RESET => n15, Q => 
                           Q(106));
   D_I_107 : FD_1362 port map( D => d(107), CK => n43, RESET => n15, Q => 
                           Q(107));
   D_I_108 : FD_1361 port map( D => d(108), CK => n43, RESET => n16, Q => 
                           Q(108));
   D_I_109 : FD_1360 port map( D => d(109), CK => n43, RESET => n16, Q => 
                           Q(109));
   D_I_110 : FD_1359 port map( D => d(110), CK => n44, RESET => n16, Q => 
                           Q(110));
   D_I_111 : FD_1358 port map( D => d(111), CK => n44, RESET => n16, Q => 
                           Q(111));
   D_I_112 : FD_1357 port map( D => d(112), CK => n44, RESET => n16, Q => 
                           Q(112));
   D_I_113 : FD_1356 port map( D => d(113), CK => n44, RESET => n16, Q => 
                           Q(113));
   D_I_114 : FD_1355 port map( D => d(114), CK => n44, RESET => n16, Q => 
                           Q(114));
   D_I_115 : FD_1354 port map( D => d(115), CK => n44, RESET => n16, Q => 
                           Q(115));
   D_I_116 : FD_1353 port map( D => d(116), CK => n44, RESET => n16, Q => 
                           Q(116));
   D_I_117 : FD_1352 port map( D => d(117), CK => n44, RESET => n16, Q => 
                           Q(117));
   D_I_118 : FD_1351 port map( D => d(118), CK => n44, RESET => n16, Q => 
                           Q(118));
   D_I_119 : FD_1350 port map( D => d(119), CK => n44, RESET => n16, Q => 
                           Q(119));
   D_I_120 : FD_1349 port map( D => d(120), CK => n44, RESET => n17, Q => 
                           Q(120));
   D_I_121 : FD_1348 port map( D => d(121), CK => n45, RESET => n17, Q => 
                           Q(121));
   D_I_122 : FD_1347 port map( D => d(122), CK => n45, RESET => n17, Q => 
                           Q(122));
   D_I_123 : FD_1346 port map( D => d(123), CK => n45, RESET => n17, Q => 
                           Q(123));
   D_I_124 : FD_1345 port map( D => d(124), CK => n45, RESET => n17, Q => 
                           Q(124));
   D_I_125 : FD_1344 port map( D => d(125), CK => n45, RESET => n17, Q => 
                           Q(125));
   D_I_126 : FD_1343 port map( D => d(126), CK => n45, RESET => n17, Q => 
                           Q(126));
   D_I_127 : FD_1342 port map( D => d(127), CK => n45, RESET => n17, Q => 
                           Q(127));
   D_I_128 : FD_1341 port map( D => d(128), CK => n45, RESET => n17, Q => 
                           Q(128));
   D_I_129 : FD_1340 port map( D => d(129), CK => n45, RESET => n17, Q => 
                           Q(129));
   D_I_130 : FD_1339 port map( D => d(130), CK => n45, RESET => n17, Q => 
                           Q(130));
   D_I_131 : FD_1338 port map( D => d(131), CK => n45, RESET => n17, Q => 
                           Q(131));
   D_I_132 : FD_1337 port map( D => d(132), CK => n46, RESET => n18, Q => 
                           Q(132));
   D_I_133 : FD_1336 port map( D => d(133), CK => n46, RESET => n18, Q => 
                           Q(133));
   D_I_134 : FD_1335 port map( D => d(134), CK => n46, RESET => n18, Q => 
                           Q(134));
   D_I_135 : FD_1334 port map( D => d(135), CK => n46, RESET => n18, Q => 
                           Q(135));
   D_I_136 : FD_1333 port map( D => d(136), CK => n46, RESET => n18, Q => 
                           Q(136));
   D_I_137 : FD_1332 port map( D => d(137), CK => n46, RESET => n18, Q => 
                           Q(137));
   D_I_138 : FD_1331 port map( D => d(138), CK => n46, RESET => n18, Q => 
                           Q(138));
   D_I_139 : FD_1330 port map( D => d(139), CK => n46, RESET => n18, Q => 
                           Q(139));
   D_I_140 : FD_1329 port map( D => d(140), CK => n46, RESET => n18, Q => 
                           Q(140));
   D_I_141 : FD_1328 port map( D => d(141), CK => n46, RESET => n18, Q => 
                           Q(141));
   D_I_142 : FD_1327 port map( D => d(142), CK => n46, RESET => n18, Q => 
                           Q(142));
   D_I_143 : FD_1326 port map( D => d(143), CK => n47, RESET => n18, Q => 
                           Q(143));
   D_I_144 : FD_1325 port map( D => d(144), CK => n47, RESET => n19, Q => 
                           Q(144));
   D_I_145 : FD_1324 port map( D => d(145), CK => n47, RESET => n19, Q => 
                           Q(145));
   D_I_146 : FD_1323 port map( D => d(146), CK => n47, RESET => n19, Q => 
                           Q(146));
   D_I_147 : FD_1322 port map( D => d(147), CK => n47, RESET => n19, Q => 
                           Q(147));
   D_I_148 : FD_1321 port map( D => d(148), CK => n47, RESET => n19, Q => 
                           Q(148));
   D_I_149 : FD_1320 port map( D => d(149), CK => n47, RESET => n19, Q => 
                           Q(149));
   D_I_150 : FD_1319 port map( D => d(150), CK => n47, RESET => n19, Q => 
                           Q(150));
   D_I_151 : FD_1318 port map( D => d(151), CK => n47, RESET => n19, Q => 
                           Q(151));
   D_I_152 : FD_1317 port map( D => d(152), CK => n47, RESET => n19, Q => 
                           Q(152));
   D_I_153 : FD_1316 port map( D => d(153), CK => n47, RESET => n19, Q => 
                           Q(153));
   D_I_154 : FD_1315 port map( D => d(154), CK => n48, RESET => n19, Q => 
                           Q(154));
   D_I_155 : FD_1314 port map( D => d(155), CK => n48, RESET => n19, Q => 
                           Q(155));
   D_I_156 : FD_1313 port map( D => d(156), CK => n48, RESET => n20, Q => 
                           Q(156));
   D_I_157 : FD_1312 port map( D => d(157), CK => n48, RESET => n20, Q => 
                           Q(157));
   D_I_158 : FD_1311 port map( D => d(158), CK => n48, RESET => n20, Q => 
                           Q(158));
   D_I_159 : FD_1310 port map( D => d(159), CK => n48, RESET => n20, Q => 
                           Q(159));
   D_I_160 : FD_1309 port map( D => d(160), CK => n48, RESET => n20, Q => 
                           Q(160));
   D_I_161 : FD_1308 port map( D => d(161), CK => n48, RESET => n20, Q => 
                           Q(161));
   D_I_162 : FD_1307 port map( D => d(162), CK => n48, RESET => n20, Q => 
                           Q(162));
   D_I_163 : FD_1306 port map( D => d(163), CK => n48, RESET => n20, Q => 
                           Q(163));
   D_I_164 : FD_1305 port map( D => d(164), CK => n48, RESET => n20, Q => 
                           Q(164));
   D_I_165 : FD_1304 port map( D => d(165), CK => n49, RESET => n20, Q => 
                           Q(165));
   D_I_166 : FD_1303 port map( D => d(166), CK => n49, RESET => n20, Q => 
                           Q(166));
   D_I_167 : FD_1302 port map( D => d(167), CK => n49, RESET => n20, Q => 
                           Q(167));
   D_I_168 : FD_1301 port map( D => d(168), CK => n49, RESET => n21, Q => 
                           Q(168));
   D_I_169 : FD_1300 port map( D => d(169), CK => n49, RESET => n21, Q => 
                           Q(169));
   D_I_170 : FD_1299 port map( D => d(170), CK => n49, RESET => n21, Q => 
                           Q(170));
   D_I_171 : FD_1298 port map( D => d(171), CK => n49, RESET => n21, Q => 
                           Q(171));
   D_I_172 : FD_1297 port map( D => d(172), CK => n49, RESET => n21, Q => 
                           Q(172));
   D_I_173 : FD_1296 port map( D => d(173), CK => n49, RESET => n21, Q => 
                           Q(173));
   D_I_174 : FD_1295 port map( D => d(174), CK => n49, RESET => n21, Q => 
                           Q(174));
   D_I_175 : FD_1294 port map( D => d(175), CK => n49, RESET => n21, Q => 
                           Q(175));
   D_I_176 : FD_1293 port map( D => d(176), CK => n50, RESET => n21, Q => 
                           Q(176));
   D_I_177 : FD_1292 port map( D => d(177), CK => n50, RESET => n21, Q => 
                           Q(177));
   D_I_178 : FD_1291 port map( D => d(178), CK => n50, RESET => n21, Q => 
                           Q(178));
   D_I_179 : FD_1290 port map( D => d(179), CK => n50, RESET => n21, Q => 
                           Q(179));
   D_I_180 : FD_1289 port map( D => d(180), CK => n50, RESET => n22, Q => 
                           Q(180));
   D_I_181 : FD_1288 port map( D => d(181), CK => n50, RESET => n22, Q => 
                           Q(181));
   D_I_182 : FD_1287 port map( D => d(182), CK => n50, RESET => n22, Q => 
                           Q(182));
   D_I_183 : FD_1286 port map( D => d(183), CK => n50, RESET => n22, Q => 
                           Q(183));
   D_I_184 : FD_1285 port map( D => d(184), CK => n50, RESET => n22, Q => 
                           Q(184));
   D_I_185 : FD_1284 port map( D => d(185), CK => n50, RESET => n22, Q => 
                           Q(185));
   D_I_186 : FD_1283 port map( D => d(186), CK => n50, RESET => n22, Q => 
                           Q(186));
   D_I_187 : FD_1282 port map( D => d(187), CK => n51, RESET => n22, Q => 
                           Q(187));
   D_I_188 : FD_1281 port map( D => d(188), CK => n51, RESET => n22, Q => 
                           Q(188));
   D_I_189 : FD_1280 port map( D => d(189), CK => n51, RESET => n22, Q => 
                           Q(189));
   D_I_190 : FD_1279 port map( D => d(190), CK => n51, RESET => n22, Q => 
                           Q(190));
   D_I_191 : FD_1278 port map( D => d(191), CK => n51, RESET => n22, Q => 
                           Q(191));
   D_I_192 : FD_1277 port map( D => d(192), CK => n51, RESET => n23, Q => 
                           Q(192));
   D_I_193 : FD_1276 port map( D => d(193), CK => n51, RESET => n23, Q => 
                           Q(193));
   D_I_194 : FD_1275 port map( D => d(194), CK => n51, RESET => n23, Q => 
                           Q(194));
   D_I_195 : FD_1274 port map( D => d(195), CK => n51, RESET => n23, Q => 
                           Q(195));
   D_I_196 : FD_1273 port map( D => d(196), CK => n51, RESET => n23, Q => 
                           Q(196));
   D_I_197 : FD_1272 port map( D => d(197), CK => n51, RESET => n23, Q => 
                           Q(197));
   D_I_198 : FD_1271 port map( D => d(198), CK => n52, RESET => n23, Q => 
                           Q(198));
   D_I_199 : FD_1270 port map( D => d(199), CK => n52, RESET => n23, Q => 
                           Q(199));
   D_I_200 : FD_1269 port map( D => d(200), CK => n52, RESET => n23, Q => 
                           Q(200));
   D_I_201 : FD_1268 port map( D => d(201), CK => n52, RESET => n23, Q => 
                           Q(201));
   D_I_202 : FD_1267 port map( D => d(202), CK => n52, RESET => n23, Q => 
                           Q(202));
   D_I_203 : FD_1266 port map( D => d(203), CK => n52, RESET => n23, Q => 
                           Q(203));
   D_I_204 : FD_1265 port map( D => d(204), CK => n52, RESET => n24, Q => 
                           Q(204));
   D_I_205 : FD_1264 port map( D => d(205), CK => n52, RESET => n24, Q => 
                           Q(205));
   D_I_206 : FD_1263 port map( D => d(206), CK => n52, RESET => n24, Q => 
                           Q(206));
   D_I_207 : FD_1262 port map( D => d(207), CK => n52, RESET => n24, Q => 
                           Q(207));
   D_I_208 : FD_1261 port map( D => d(208), CK => n52, RESET => n24, Q => 
                           Q(208));
   D_I_209 : FD_1260 port map( D => d(209), CK => n53, RESET => n24, Q => 
                           Q(209));
   D_I_210 : FD_1259 port map( D => d(210), CK => n53, RESET => n24, Q => 
                           Q(210));
   D_I_211 : FD_1258 port map( D => d(211), CK => n53, RESET => n24, Q => 
                           Q(211));
   D_I_212 : FD_1257 port map( D => d(212), CK => n53, RESET => n24, Q => 
                           Q(212));
   D_I_213 : FD_1256 port map( D => d(213), CK => n53, RESET => n24, Q => 
                           Q(213));
   D_I_214 : FD_1255 port map( D => d(214), CK => n53, RESET => n24, Q => 
                           Q(214));
   D_I_215 : FD_1254 port map( D => d(215), CK => n53, RESET => n24, Q => 
                           Q(215));
   D_I_216 : FD_1253 port map( D => d(216), CK => n53, RESET => n25, Q => 
                           Q(216));
   D_I_217 : FD_1252 port map( D => d(217), CK => n53, RESET => n25, Q => 
                           Q(217));
   D_I_218 : FD_1251 port map( D => d(218), CK => n53, RESET => n25, Q => 
                           Q(218));
   D_I_219 : FD_1250 port map( D => d(219), CK => n53, RESET => n25, Q => 
                           Q(219));
   D_I_220 : FD_1249 port map( D => d(220), CK => n54, RESET => n25, Q => 
                           Q(220));
   D_I_221 : FD_1248 port map( D => d(221), CK => n54, RESET => n25, Q => 
                           Q(221));
   D_I_222 : FD_1247 port map( D => d(222), CK => n54, RESET => n25, Q => 
                           Q(222));
   D_I_223 : FD_1246 port map( D => d(223), CK => n54, RESET => n25, Q => 
                           Q(223));
   D_I_224 : FD_1245 port map( D => d(224), CK => n54, RESET => n25, Q => 
                           Q(224));
   D_I_225 : FD_1244 port map( D => d(225), CK => n54, RESET => n25, Q => 
                           Q(225));
   D_I_226 : FD_1243 port map( D => d(226), CK => n54, RESET => n25, Q => 
                           Q(226));
   D_I_227 : FD_1242 port map( D => d(227), CK => n54, RESET => n25, Q => 
                           Q(227));
   D_I_228 : FD_1241 port map( D => d(228), CK => n54, RESET => n26, Q => 
                           Q(228));
   D_I_229 : FD_1240 port map( D => d(229), CK => n54, RESET => n26, Q => 
                           Q(229));
   D_I_230 : FD_1239 port map( D => d(230), CK => n54, RESET => n26, Q => 
                           Q(230));
   D_I_231 : FD_1238 port map( D => d(231), CK => n55, RESET => n26, Q => 
                           Q(231));
   D_I_232 : FD_1237 port map( D => d(232), CK => n55, RESET => n26, Q => 
                           Q(232));
   D_I_233 : FD_1236 port map( D => d(233), CK => n55, RESET => n26, Q => 
                           Q(233));
   D_I_234 : FD_1235 port map( D => d(234), CK => n55, RESET => n26, Q => 
                           Q(234));
   D_I_235 : FD_1234 port map( D => d(235), CK => n55, RESET => n26, Q => 
                           Q(235));
   D_I_236 : FD_1233 port map( D => d(236), CK => n55, RESET => n26, Q => 
                           Q(236));
   D_I_237 : FD_1232 port map( D => d(237), CK => n55, RESET => n26, Q => 
                           Q(237));
   D_I_238 : FD_1231 port map( D => d(238), CK => n55, RESET => n26, Q => 
                           Q(238));
   D_I_239 : FD_1230 port map( D => d(239), CK => n55, RESET => n26, Q => 
                           Q(239));
   D_I_240 : FD_1229 port map( D => d(240), CK => n55, RESET => n27, Q => 
                           Q(240));
   D_I_241 : FD_1228 port map( D => d(241), CK => n55, RESET => n27, Q => 
                           Q(241));
   D_I_242 : FD_1227 port map( D => d(242), CK => n56, RESET => n27, Q => 
                           Q(242));
   D_I_243 : FD_1226 port map( D => d(243), CK => n56, RESET => n27, Q => 
                           Q(243));
   D_I_244 : FD_1225 port map( D => d(244), CK => n56, RESET => n27, Q => 
                           Q(244));
   D_I_245 : FD_1224 port map( D => d(245), CK => n56, RESET => n27, Q => 
                           Q(245));
   D_I_246 : FD_1223 port map( D => d(246), CK => n56, RESET => n27, Q => 
                           Q(246));
   D_I_247 : FD_1222 port map( D => d(247), CK => n56, RESET => n27, Q => 
                           Q(247));
   D_I_248 : FD_1221 port map( D => d(248), CK => n56, RESET => n27, Q => 
                           Q(248));
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_4 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_4;

architecture SYN_struc of reg_nbit_n249_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_940
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_941
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_942
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_943
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_944
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_945
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_946
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_947
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_948
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_949
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_950
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_951
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_952
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_953
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_954
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_955
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_956
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_957
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_958
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_959
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_960
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_961
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_962
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_963
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_964
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_965
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_966
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_967
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_968
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_969
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_970
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_971
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_972
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_973
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_974
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_975
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_976
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_977
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_978
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_979
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_980
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_981
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_982
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_983
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_984
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_985
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_986
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_987
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_988
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_989
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_990
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_991
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_992
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_993
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_994
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_995
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_996
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_997
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_998
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_999
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1000
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1001
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1002
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1003
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1004
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1005
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1006
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1007
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1008
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1009
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1010
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1011
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1012
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1013
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1014
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1015
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1016
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1017
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1018
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1019
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1020
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1021
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1022
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1023
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1024
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1025
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1026
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1027
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1028
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1029
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1030
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1031
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1032
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1033
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1034
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1035
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1036
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1037
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1038
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1039
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1040
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1041
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1042
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1043
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1044
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1045
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1046
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1047
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1048
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1049
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1050
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1051
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1052
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1053
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1054
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1055
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1056
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1057
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1058
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1059
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1060
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1061
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1062
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1063
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1064
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1065
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1066
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1067
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1068
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1069
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1070
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1071
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1072
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1073
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1074
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1075
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1076
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1077
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1078
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1079
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1080
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1081
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1082
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1083
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1084
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1085
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1086
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1087
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1088
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1089
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1090
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1091
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1092
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1093
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1094
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1095
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1096
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1097
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1098
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1099
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1100
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1101
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1102
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1103
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1104
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1105
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1106
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1107
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1108
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1109
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1110
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1111
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1112
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1113
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1114
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1115
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1116
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1117
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1118
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1119
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1120
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1121
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1122
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1123
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1124
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1125
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1126
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1127
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1128
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1129
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1130
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1131
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1132
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1133
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1134
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1135
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1136
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1137
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1138
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1139
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1140
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1141
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1142
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1143
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1144
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1145
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1146
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1147
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1148
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1149
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1150
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1151
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1152
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1153
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1154
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1155
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1156
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1157
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1158
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1159
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1160
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1161
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1162
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1163
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1164
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1165
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1166
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1167
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1168
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1169
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1170
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1171
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1172
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1173
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1174
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1175
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1176
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1177
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1178
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1179
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1180
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1181
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1182
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1183
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1184
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1185
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1186
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1187
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1188
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_1188 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_1187 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_1186 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_1185 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_1184 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_1183 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_1182 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_1181 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_1180 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_1179 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_1178 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_1177 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_1176 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_1175 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_1174 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_1173 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_1172 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_1171 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_1170 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_1169 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_1168 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_1167 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_1166 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_1165 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_1164 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_1163 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_1162 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_1161 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_1160 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_1159 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_1158 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_1157 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_1156 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_1155 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_1154 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_1153 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_1152 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_1151 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_1150 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_1149 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_1148 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_1147 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_1146 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_1145 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_1144 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_1143 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_1142 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_1141 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_1140 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_1139 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_1138 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_1137 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_1136 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_1135 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_1134 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_1133 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_1132 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_1131 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_1130 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_1129 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_1128 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_1127 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_1126 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_1125 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_1124 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_1123 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_1122 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_1121 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_1120 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_1119 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_1118 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_1117 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_1116 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_1115 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_1114 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_1113 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_1112 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_1111 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_1110 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_1109 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_1108 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_1107 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_1106 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_1105 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_1104 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_1103 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_1102 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_1101 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_1100 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_1099 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_1098 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_1097 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_1096 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_1095 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_1094 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_1093 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_1092 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_1091 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_1090 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_1089 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_1088 port map( D => d(100), CK => n43, RESET => n15, Q => 
                           Q(100));
   D_I_101 : FD_1087 port map( D => d(101), CK => n43, RESET => n15, Q => 
                           Q(101));
   D_I_102 : FD_1086 port map( D => d(102), CK => n43, RESET => n15, Q => 
                           Q(102));
   D_I_103 : FD_1085 port map( D => d(103), CK => n43, RESET => n15, Q => 
                           Q(103));
   D_I_104 : FD_1084 port map( D => d(104), CK => n43, RESET => n15, Q => 
                           Q(104));
   D_I_105 : FD_1083 port map( D => d(105), CK => n43, RESET => n15, Q => 
                           Q(105));
   D_I_106 : FD_1082 port map( D => d(106), CK => n43, RESET => n15, Q => 
                           Q(106));
   D_I_107 : FD_1081 port map( D => d(107), CK => n43, RESET => n15, Q => 
                           Q(107));
   D_I_108 : FD_1080 port map( D => d(108), CK => n43, RESET => n16, Q => 
                           Q(108));
   D_I_109 : FD_1079 port map( D => d(109), CK => n43, RESET => n16, Q => 
                           Q(109));
   D_I_110 : FD_1078 port map( D => d(110), CK => n44, RESET => n16, Q => 
                           Q(110));
   D_I_111 : FD_1077 port map( D => d(111), CK => n44, RESET => n16, Q => 
                           Q(111));
   D_I_112 : FD_1076 port map( D => d(112), CK => n44, RESET => n16, Q => 
                           Q(112));
   D_I_113 : FD_1075 port map( D => d(113), CK => n44, RESET => n16, Q => 
                           Q(113));
   D_I_114 : FD_1074 port map( D => d(114), CK => n44, RESET => n16, Q => 
                           Q(114));
   D_I_115 : FD_1073 port map( D => d(115), CK => n44, RESET => n16, Q => 
                           Q(115));
   D_I_116 : FD_1072 port map( D => d(116), CK => n44, RESET => n16, Q => 
                           Q(116));
   D_I_117 : FD_1071 port map( D => d(117), CK => n44, RESET => n16, Q => 
                           Q(117));
   D_I_118 : FD_1070 port map( D => d(118), CK => n44, RESET => n16, Q => 
                           Q(118));
   D_I_119 : FD_1069 port map( D => d(119), CK => n44, RESET => n16, Q => 
                           Q(119));
   D_I_120 : FD_1068 port map( D => d(120), CK => n44, RESET => n17, Q => 
                           Q(120));
   D_I_121 : FD_1067 port map( D => d(121), CK => n45, RESET => n17, Q => 
                           Q(121));
   D_I_122 : FD_1066 port map( D => d(122), CK => n45, RESET => n17, Q => 
                           Q(122));
   D_I_123 : FD_1065 port map( D => d(123), CK => n45, RESET => n17, Q => 
                           Q(123));
   D_I_124 : FD_1064 port map( D => d(124), CK => n45, RESET => n17, Q => 
                           Q(124));
   D_I_125 : FD_1063 port map( D => d(125), CK => n45, RESET => n17, Q => 
                           Q(125));
   D_I_126 : FD_1062 port map( D => d(126), CK => n45, RESET => n17, Q => 
                           Q(126));
   D_I_127 : FD_1061 port map( D => d(127), CK => n45, RESET => n17, Q => 
                           Q(127));
   D_I_128 : FD_1060 port map( D => d(128), CK => n45, RESET => n17, Q => 
                           Q(128));
   D_I_129 : FD_1059 port map( D => d(129), CK => n45, RESET => n17, Q => 
                           Q(129));
   D_I_130 : FD_1058 port map( D => d(130), CK => n45, RESET => n17, Q => 
                           Q(130));
   D_I_131 : FD_1057 port map( D => d(131), CK => n45, RESET => n17, Q => 
                           Q(131));
   D_I_132 : FD_1056 port map( D => d(132), CK => n46, RESET => n18, Q => 
                           Q(132));
   D_I_133 : FD_1055 port map( D => d(133), CK => n46, RESET => n18, Q => 
                           Q(133));
   D_I_134 : FD_1054 port map( D => d(134), CK => n46, RESET => n18, Q => 
                           Q(134));
   D_I_135 : FD_1053 port map( D => d(135), CK => n46, RESET => n18, Q => 
                           Q(135));
   D_I_136 : FD_1052 port map( D => d(136), CK => n46, RESET => n18, Q => 
                           Q(136));
   D_I_137 : FD_1051 port map( D => d(137), CK => n46, RESET => n18, Q => 
                           Q(137));
   D_I_138 : FD_1050 port map( D => d(138), CK => n46, RESET => n18, Q => 
                           Q(138));
   D_I_139 : FD_1049 port map( D => d(139), CK => n46, RESET => n18, Q => 
                           Q(139));
   D_I_140 : FD_1048 port map( D => d(140), CK => n46, RESET => n18, Q => 
                           Q(140));
   D_I_141 : FD_1047 port map( D => d(141), CK => n46, RESET => n18, Q => 
                           Q(141));
   D_I_142 : FD_1046 port map( D => d(142), CK => n46, RESET => n18, Q => 
                           Q(142));
   D_I_143 : FD_1045 port map( D => d(143), CK => n47, RESET => n18, Q => 
                           Q(143));
   D_I_144 : FD_1044 port map( D => d(144), CK => n47, RESET => n19, Q => 
                           Q(144));
   D_I_145 : FD_1043 port map( D => d(145), CK => n47, RESET => n19, Q => 
                           Q(145));
   D_I_146 : FD_1042 port map( D => d(146), CK => n47, RESET => n19, Q => 
                           Q(146));
   D_I_147 : FD_1041 port map( D => d(147), CK => n47, RESET => n19, Q => 
                           Q(147));
   D_I_148 : FD_1040 port map( D => d(148), CK => n47, RESET => n19, Q => 
                           Q(148));
   D_I_149 : FD_1039 port map( D => d(149), CK => n47, RESET => n19, Q => 
                           Q(149));
   D_I_150 : FD_1038 port map( D => d(150), CK => n47, RESET => n19, Q => 
                           Q(150));
   D_I_151 : FD_1037 port map( D => d(151), CK => n47, RESET => n19, Q => 
                           Q(151));
   D_I_152 : FD_1036 port map( D => d(152), CK => n47, RESET => n19, Q => 
                           Q(152));
   D_I_153 : FD_1035 port map( D => d(153), CK => n47, RESET => n19, Q => 
                           Q(153));
   D_I_154 : FD_1034 port map( D => d(154), CK => n48, RESET => n19, Q => 
                           Q(154));
   D_I_155 : FD_1033 port map( D => d(155), CK => n48, RESET => n19, Q => 
                           Q(155));
   D_I_156 : FD_1032 port map( D => d(156), CK => n48, RESET => n20, Q => 
                           Q(156));
   D_I_157 : FD_1031 port map( D => d(157), CK => n48, RESET => n20, Q => 
                           Q(157));
   D_I_158 : FD_1030 port map( D => d(158), CK => n48, RESET => n20, Q => 
                           Q(158));
   D_I_159 : FD_1029 port map( D => d(159), CK => n48, RESET => n20, Q => 
                           Q(159));
   D_I_160 : FD_1028 port map( D => d(160), CK => n48, RESET => n20, Q => 
                           Q(160));
   D_I_161 : FD_1027 port map( D => d(161), CK => n48, RESET => n20, Q => 
                           Q(161));
   D_I_162 : FD_1026 port map( D => d(162), CK => n48, RESET => n20, Q => 
                           Q(162));
   D_I_163 : FD_1025 port map( D => d(163), CK => n48, RESET => n20, Q => 
                           Q(163));
   D_I_164 : FD_1024 port map( D => d(164), CK => n48, RESET => n20, Q => 
                           Q(164));
   D_I_165 : FD_1023 port map( D => d(165), CK => n49, RESET => n20, Q => 
                           Q(165));
   D_I_166 : FD_1022 port map( D => d(166), CK => n49, RESET => n20, Q => 
                           Q(166));
   D_I_167 : FD_1021 port map( D => d(167), CK => n49, RESET => n20, Q => 
                           Q(167));
   D_I_168 : FD_1020 port map( D => d(168), CK => n49, RESET => n21, Q => 
                           Q(168));
   D_I_169 : FD_1019 port map( D => d(169), CK => n49, RESET => n21, Q => 
                           Q(169));
   D_I_170 : FD_1018 port map( D => d(170), CK => n49, RESET => n21, Q => 
                           Q(170));
   D_I_171 : FD_1017 port map( D => d(171), CK => n49, RESET => n21, Q => 
                           Q(171));
   D_I_172 : FD_1016 port map( D => d(172), CK => n49, RESET => n21, Q => 
                           Q(172));
   D_I_173 : FD_1015 port map( D => d(173), CK => n49, RESET => n21, Q => 
                           Q(173));
   D_I_174 : FD_1014 port map( D => d(174), CK => n49, RESET => n21, Q => 
                           Q(174));
   D_I_175 : FD_1013 port map( D => d(175), CK => n49, RESET => n21, Q => 
                           Q(175));
   D_I_176 : FD_1012 port map( D => d(176), CK => n50, RESET => n21, Q => 
                           Q(176));
   D_I_177 : FD_1011 port map( D => d(177), CK => n50, RESET => n21, Q => 
                           Q(177));
   D_I_178 : FD_1010 port map( D => d(178), CK => n50, RESET => n21, Q => 
                           Q(178));
   D_I_179 : FD_1009 port map( D => d(179), CK => n50, RESET => n21, Q => 
                           Q(179));
   D_I_180 : FD_1008 port map( D => d(180), CK => n50, RESET => n22, Q => 
                           Q(180));
   D_I_181 : FD_1007 port map( D => d(181), CK => n50, RESET => n22, Q => 
                           Q(181));
   D_I_182 : FD_1006 port map( D => d(182), CK => n50, RESET => n22, Q => 
                           Q(182));
   D_I_183 : FD_1005 port map( D => d(183), CK => n50, RESET => n22, Q => 
                           Q(183));
   D_I_184 : FD_1004 port map( D => d(184), CK => n50, RESET => n22, Q => 
                           Q(184));
   D_I_185 : FD_1003 port map( D => d(185), CK => n50, RESET => n22, Q => 
                           Q(185));
   D_I_186 : FD_1002 port map( D => d(186), CK => n50, RESET => n22, Q => 
                           Q(186));
   D_I_187 : FD_1001 port map( D => d(187), CK => n51, RESET => n22, Q => 
                           Q(187));
   D_I_188 : FD_1000 port map( D => d(188), CK => n51, RESET => n22, Q => 
                           Q(188));
   D_I_189 : FD_999 port map( D => d(189), CK => n51, RESET => n22, Q => Q(189)
                           );
   D_I_190 : FD_998 port map( D => d(190), CK => n51, RESET => n22, Q => Q(190)
                           );
   D_I_191 : FD_997 port map( D => d(191), CK => n51, RESET => n22, Q => Q(191)
                           );
   D_I_192 : FD_996 port map( D => d(192), CK => n51, RESET => n23, Q => Q(192)
                           );
   D_I_193 : FD_995 port map( D => d(193), CK => n51, RESET => n23, Q => Q(193)
                           );
   D_I_194 : FD_994 port map( D => d(194), CK => n51, RESET => n23, Q => Q(194)
                           );
   D_I_195 : FD_993 port map( D => d(195), CK => n51, RESET => n23, Q => Q(195)
                           );
   D_I_196 : FD_992 port map( D => d(196), CK => n51, RESET => n23, Q => Q(196)
                           );
   D_I_197 : FD_991 port map( D => d(197), CK => n51, RESET => n23, Q => Q(197)
                           );
   D_I_198 : FD_990 port map( D => d(198), CK => n52, RESET => n23, Q => Q(198)
                           );
   D_I_199 : FD_989 port map( D => d(199), CK => n52, RESET => n23, Q => Q(199)
                           );
   D_I_200 : FD_988 port map( D => d(200), CK => n52, RESET => n23, Q => Q(200)
                           );
   D_I_201 : FD_987 port map( D => d(201), CK => n52, RESET => n23, Q => Q(201)
                           );
   D_I_202 : FD_986 port map( D => d(202), CK => n52, RESET => n23, Q => Q(202)
                           );
   D_I_203 : FD_985 port map( D => d(203), CK => n52, RESET => n23, Q => Q(203)
                           );
   D_I_204 : FD_984 port map( D => d(204), CK => n52, RESET => n24, Q => Q(204)
                           );
   D_I_205 : FD_983 port map( D => d(205), CK => n52, RESET => n24, Q => Q(205)
                           );
   D_I_206 : FD_982 port map( D => d(206), CK => n52, RESET => n24, Q => Q(206)
                           );
   D_I_207 : FD_981 port map( D => d(207), CK => n52, RESET => n24, Q => Q(207)
                           );
   D_I_208 : FD_980 port map( D => d(208), CK => n52, RESET => n24, Q => Q(208)
                           );
   D_I_209 : FD_979 port map( D => d(209), CK => n53, RESET => n24, Q => Q(209)
                           );
   D_I_210 : FD_978 port map( D => d(210), CK => n53, RESET => n24, Q => Q(210)
                           );
   D_I_211 : FD_977 port map( D => d(211), CK => n53, RESET => n24, Q => Q(211)
                           );
   D_I_212 : FD_976 port map( D => d(212), CK => n53, RESET => n24, Q => Q(212)
                           );
   D_I_213 : FD_975 port map( D => d(213), CK => n53, RESET => n24, Q => Q(213)
                           );
   D_I_214 : FD_974 port map( D => d(214), CK => n53, RESET => n24, Q => Q(214)
                           );
   D_I_215 : FD_973 port map( D => d(215), CK => n53, RESET => n24, Q => Q(215)
                           );
   D_I_216 : FD_972 port map( D => d(216), CK => n53, RESET => n25, Q => Q(216)
                           );
   D_I_217 : FD_971 port map( D => d(217), CK => n53, RESET => n25, Q => Q(217)
                           );
   D_I_218 : FD_970 port map( D => d(218), CK => n53, RESET => n25, Q => Q(218)
                           );
   D_I_219 : FD_969 port map( D => d(219), CK => n53, RESET => n25, Q => Q(219)
                           );
   D_I_220 : FD_968 port map( D => d(220), CK => n54, RESET => n25, Q => Q(220)
                           );
   D_I_221 : FD_967 port map( D => d(221), CK => n54, RESET => n25, Q => Q(221)
                           );
   D_I_222 : FD_966 port map( D => d(222), CK => n54, RESET => n25, Q => Q(222)
                           );
   D_I_223 : FD_965 port map( D => d(223), CK => n54, RESET => n25, Q => Q(223)
                           );
   D_I_224 : FD_964 port map( D => d(224), CK => n54, RESET => n25, Q => Q(224)
                           );
   D_I_225 : FD_963 port map( D => d(225), CK => n54, RESET => n25, Q => Q(225)
                           );
   D_I_226 : FD_962 port map( D => d(226), CK => n54, RESET => n25, Q => Q(226)
                           );
   D_I_227 : FD_961 port map( D => d(227), CK => n54, RESET => n25, Q => Q(227)
                           );
   D_I_228 : FD_960 port map( D => d(228), CK => n54, RESET => n26, Q => Q(228)
                           );
   D_I_229 : FD_959 port map( D => d(229), CK => n54, RESET => n26, Q => Q(229)
                           );
   D_I_230 : FD_958 port map( D => d(230), CK => n54, RESET => n26, Q => Q(230)
                           );
   D_I_231 : FD_957 port map( D => d(231), CK => n55, RESET => n26, Q => Q(231)
                           );
   D_I_232 : FD_956 port map( D => d(232), CK => n55, RESET => n26, Q => Q(232)
                           );
   D_I_233 : FD_955 port map( D => d(233), CK => n55, RESET => n26, Q => Q(233)
                           );
   D_I_234 : FD_954 port map( D => d(234), CK => n55, RESET => n26, Q => Q(234)
                           );
   D_I_235 : FD_953 port map( D => d(235), CK => n55, RESET => n26, Q => Q(235)
                           );
   D_I_236 : FD_952 port map( D => d(236), CK => n55, RESET => n26, Q => Q(236)
                           );
   D_I_237 : FD_951 port map( D => d(237), CK => n55, RESET => n26, Q => Q(237)
                           );
   D_I_238 : FD_950 port map( D => d(238), CK => n55, RESET => n26, Q => Q(238)
                           );
   D_I_239 : FD_949 port map( D => d(239), CK => n55, RESET => n26, Q => Q(239)
                           );
   D_I_240 : FD_948 port map( D => d(240), CK => n55, RESET => n27, Q => Q(240)
                           );
   D_I_241 : FD_947 port map( D => d(241), CK => n55, RESET => n27, Q => Q(241)
                           );
   D_I_242 : FD_946 port map( D => d(242), CK => n56, RESET => n27, Q => Q(242)
                           );
   D_I_243 : FD_945 port map( D => d(243), CK => n56, RESET => n27, Q => Q(243)
                           );
   D_I_244 : FD_944 port map( D => d(244), CK => n56, RESET => n27, Q => Q(244)
                           );
   D_I_245 : FD_943 port map( D => d(245), CK => n56, RESET => n27, Q => Q(245)
                           );
   D_I_246 : FD_942 port map( D => d(246), CK => n56, RESET => n27, Q => Q(246)
                           );
   D_I_247 : FD_941 port map( D => d(247), CK => n56, RESET => n27, Q => Q(247)
                           );
   D_I_248 : FD_940 port map( D => d(248), CK => n56, RESET => n27, Q => Q(248)
                           );
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_3 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_3;

architecture SYN_struc of reg_nbit_n249_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_659
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_660
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_661
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_662
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_663
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_664
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_665
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_666
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_667
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_668
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_669
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_670
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_671
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_672
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_673
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_674
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_675
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_676
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_677
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_678
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_679
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_680
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_681
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_682
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_683
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_684
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_685
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_686
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_687
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_688
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_689
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_690
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_691
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_692
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_693
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_694
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_695
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_696
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_697
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_698
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_699
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_700
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_701
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_702
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_703
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_704
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_705
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_706
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_707
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_708
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_709
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_710
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_711
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_712
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_713
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_714
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_715
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_716
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_717
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_718
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_719
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_720
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_721
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_722
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_723
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_724
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_725
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_726
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_727
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_728
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_729
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_730
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_731
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_732
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_733
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_734
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_735
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_736
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_737
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_738
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_739
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_740
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_741
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_742
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_743
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_744
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_745
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_746
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_747
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_748
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_749
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_750
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_751
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_752
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_753
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_754
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_755
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_756
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_757
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_758
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_759
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_760
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_761
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_762
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_763
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_764
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_765
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_766
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_767
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_768
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_769
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_770
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_771
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_772
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_773
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_774
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_775
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_776
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_777
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_778
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_779
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_780
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_781
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_782
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_783
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_784
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_785
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_786
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_787
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_788
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_789
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_790
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_791
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_792
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_793
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_794
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_795
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_796
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_797
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_798
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_799
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_800
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_801
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_802
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_803
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_804
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_805
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_806
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_807
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_808
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_809
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_810
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_811
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_812
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_813
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_814
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_815
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_816
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_817
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_818
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_819
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_820
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_821
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_822
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_823
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_824
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_825
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_826
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_827
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_828
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_829
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_830
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_831
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_832
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_833
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_834
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_835
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_836
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_837
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_838
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_839
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_840
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_841
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_842
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_843
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_844
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_845
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_846
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_847
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_848
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_849
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_850
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_851
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_852
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_853
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_854
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_855
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_856
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_857
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_858
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_859
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_860
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_861
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_862
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_863
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_864
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_865
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_866
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_867
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_868
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_869
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_870
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_871
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_872
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_873
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_874
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_875
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_876
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_877
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_878
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_879
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_880
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_881
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_882
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_883
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_884
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_885
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_886
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_887
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_888
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_889
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_890
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_891
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_892
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_893
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_894
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_895
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_896
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_897
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_898
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_899
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_900
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_901
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_902
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_903
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_904
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_905
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_906
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_907
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_907 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_906 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_905 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_904 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_903 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_902 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_901 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_900 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_899 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_898 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_897 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_896 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_895 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_894 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_893 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_892 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_891 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_890 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_889 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_888 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_887 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_886 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_885 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_884 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_883 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_882 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_881 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_880 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_879 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_878 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_877 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_876 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_875 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_874 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_873 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_872 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_871 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_870 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_869 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_868 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_867 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_866 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_865 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_864 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_863 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_862 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_861 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_860 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_859 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_858 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_857 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_856 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_855 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_854 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_853 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_852 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_851 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_850 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_849 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_848 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_847 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_846 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_845 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_844 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_843 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_842 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_841 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_840 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_839 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_838 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_837 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_836 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_835 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_834 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_833 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_832 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_831 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_830 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_829 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_828 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_827 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_826 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_825 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_824 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_823 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_822 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_821 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_820 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_819 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_818 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_817 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_816 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_815 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_814 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_813 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_812 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_811 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_810 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_809 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_808 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_807 port map( D => d(100), CK => n43, RESET => n15, Q => Q(100)
                           );
   D_I_101 : FD_806 port map( D => d(101), CK => n43, RESET => n15, Q => Q(101)
                           );
   D_I_102 : FD_805 port map( D => d(102), CK => n43, RESET => n15, Q => Q(102)
                           );
   D_I_103 : FD_804 port map( D => d(103), CK => n43, RESET => n15, Q => Q(103)
                           );
   D_I_104 : FD_803 port map( D => d(104), CK => n43, RESET => n15, Q => Q(104)
                           );
   D_I_105 : FD_802 port map( D => d(105), CK => n43, RESET => n15, Q => Q(105)
                           );
   D_I_106 : FD_801 port map( D => d(106), CK => n43, RESET => n15, Q => Q(106)
                           );
   D_I_107 : FD_800 port map( D => d(107), CK => n43, RESET => n15, Q => Q(107)
                           );
   D_I_108 : FD_799 port map( D => d(108), CK => n43, RESET => n16, Q => Q(108)
                           );
   D_I_109 : FD_798 port map( D => d(109), CK => n43, RESET => n16, Q => Q(109)
                           );
   D_I_110 : FD_797 port map( D => d(110), CK => n44, RESET => n16, Q => Q(110)
                           );
   D_I_111 : FD_796 port map( D => d(111), CK => n44, RESET => n16, Q => Q(111)
                           );
   D_I_112 : FD_795 port map( D => d(112), CK => n44, RESET => n16, Q => Q(112)
                           );
   D_I_113 : FD_794 port map( D => d(113), CK => n44, RESET => n16, Q => Q(113)
                           );
   D_I_114 : FD_793 port map( D => d(114), CK => n44, RESET => n16, Q => Q(114)
                           );
   D_I_115 : FD_792 port map( D => d(115), CK => n44, RESET => n16, Q => Q(115)
                           );
   D_I_116 : FD_791 port map( D => d(116), CK => n44, RESET => n16, Q => Q(116)
                           );
   D_I_117 : FD_790 port map( D => d(117), CK => n44, RESET => n16, Q => Q(117)
                           );
   D_I_118 : FD_789 port map( D => d(118), CK => n44, RESET => n16, Q => Q(118)
                           );
   D_I_119 : FD_788 port map( D => d(119), CK => n44, RESET => n16, Q => Q(119)
                           );
   D_I_120 : FD_787 port map( D => d(120), CK => n44, RESET => n17, Q => Q(120)
                           );
   D_I_121 : FD_786 port map( D => d(121), CK => n45, RESET => n17, Q => Q(121)
                           );
   D_I_122 : FD_785 port map( D => d(122), CK => n45, RESET => n17, Q => Q(122)
                           );
   D_I_123 : FD_784 port map( D => d(123), CK => n45, RESET => n17, Q => Q(123)
                           );
   D_I_124 : FD_783 port map( D => d(124), CK => n45, RESET => n17, Q => Q(124)
                           );
   D_I_125 : FD_782 port map( D => d(125), CK => n45, RESET => n17, Q => Q(125)
                           );
   D_I_126 : FD_781 port map( D => d(126), CK => n45, RESET => n17, Q => Q(126)
                           );
   D_I_127 : FD_780 port map( D => d(127), CK => n45, RESET => n17, Q => Q(127)
                           );
   D_I_128 : FD_779 port map( D => d(128), CK => n45, RESET => n17, Q => Q(128)
                           );
   D_I_129 : FD_778 port map( D => d(129), CK => n45, RESET => n17, Q => Q(129)
                           );
   D_I_130 : FD_777 port map( D => d(130), CK => n45, RESET => n17, Q => Q(130)
                           );
   D_I_131 : FD_776 port map( D => d(131), CK => n45, RESET => n17, Q => Q(131)
                           );
   D_I_132 : FD_775 port map( D => d(132), CK => n46, RESET => n18, Q => Q(132)
                           );
   D_I_133 : FD_774 port map( D => d(133), CK => n46, RESET => n18, Q => Q(133)
                           );
   D_I_134 : FD_773 port map( D => d(134), CK => n46, RESET => n18, Q => Q(134)
                           );
   D_I_135 : FD_772 port map( D => d(135), CK => n46, RESET => n18, Q => Q(135)
                           );
   D_I_136 : FD_771 port map( D => d(136), CK => n46, RESET => n18, Q => Q(136)
                           );
   D_I_137 : FD_770 port map( D => d(137), CK => n46, RESET => n18, Q => Q(137)
                           );
   D_I_138 : FD_769 port map( D => d(138), CK => n46, RESET => n18, Q => Q(138)
                           );
   D_I_139 : FD_768 port map( D => d(139), CK => n46, RESET => n18, Q => Q(139)
                           );
   D_I_140 : FD_767 port map( D => d(140), CK => n46, RESET => n18, Q => Q(140)
                           );
   D_I_141 : FD_766 port map( D => d(141), CK => n46, RESET => n18, Q => Q(141)
                           );
   D_I_142 : FD_765 port map( D => d(142), CK => n46, RESET => n18, Q => Q(142)
                           );
   D_I_143 : FD_764 port map( D => d(143), CK => n47, RESET => n18, Q => Q(143)
                           );
   D_I_144 : FD_763 port map( D => d(144), CK => n47, RESET => n19, Q => Q(144)
                           );
   D_I_145 : FD_762 port map( D => d(145), CK => n47, RESET => n19, Q => Q(145)
                           );
   D_I_146 : FD_761 port map( D => d(146), CK => n47, RESET => n19, Q => Q(146)
                           );
   D_I_147 : FD_760 port map( D => d(147), CK => n47, RESET => n19, Q => Q(147)
                           );
   D_I_148 : FD_759 port map( D => d(148), CK => n47, RESET => n19, Q => Q(148)
                           );
   D_I_149 : FD_758 port map( D => d(149), CK => n47, RESET => n19, Q => Q(149)
                           );
   D_I_150 : FD_757 port map( D => d(150), CK => n47, RESET => n19, Q => Q(150)
                           );
   D_I_151 : FD_756 port map( D => d(151), CK => n47, RESET => n19, Q => Q(151)
                           );
   D_I_152 : FD_755 port map( D => d(152), CK => n47, RESET => n19, Q => Q(152)
                           );
   D_I_153 : FD_754 port map( D => d(153), CK => n47, RESET => n19, Q => Q(153)
                           );
   D_I_154 : FD_753 port map( D => d(154), CK => n48, RESET => n19, Q => Q(154)
                           );
   D_I_155 : FD_752 port map( D => d(155), CK => n48, RESET => n19, Q => Q(155)
                           );
   D_I_156 : FD_751 port map( D => d(156), CK => n48, RESET => n20, Q => Q(156)
                           );
   D_I_157 : FD_750 port map( D => d(157), CK => n48, RESET => n20, Q => Q(157)
                           );
   D_I_158 : FD_749 port map( D => d(158), CK => n48, RESET => n20, Q => Q(158)
                           );
   D_I_159 : FD_748 port map( D => d(159), CK => n48, RESET => n20, Q => Q(159)
                           );
   D_I_160 : FD_747 port map( D => d(160), CK => n48, RESET => n20, Q => Q(160)
                           );
   D_I_161 : FD_746 port map( D => d(161), CK => n48, RESET => n20, Q => Q(161)
                           );
   D_I_162 : FD_745 port map( D => d(162), CK => n48, RESET => n20, Q => Q(162)
                           );
   D_I_163 : FD_744 port map( D => d(163), CK => n48, RESET => n20, Q => Q(163)
                           );
   D_I_164 : FD_743 port map( D => d(164), CK => n48, RESET => n20, Q => Q(164)
                           );
   D_I_165 : FD_742 port map( D => d(165), CK => n49, RESET => n20, Q => Q(165)
                           );
   D_I_166 : FD_741 port map( D => d(166), CK => n49, RESET => n20, Q => Q(166)
                           );
   D_I_167 : FD_740 port map( D => d(167), CK => n49, RESET => n20, Q => Q(167)
                           );
   D_I_168 : FD_739 port map( D => d(168), CK => n49, RESET => n21, Q => Q(168)
                           );
   D_I_169 : FD_738 port map( D => d(169), CK => n49, RESET => n21, Q => Q(169)
                           );
   D_I_170 : FD_737 port map( D => d(170), CK => n49, RESET => n21, Q => Q(170)
                           );
   D_I_171 : FD_736 port map( D => d(171), CK => n49, RESET => n21, Q => Q(171)
                           );
   D_I_172 : FD_735 port map( D => d(172), CK => n49, RESET => n21, Q => Q(172)
                           );
   D_I_173 : FD_734 port map( D => d(173), CK => n49, RESET => n21, Q => Q(173)
                           );
   D_I_174 : FD_733 port map( D => d(174), CK => n49, RESET => n21, Q => Q(174)
                           );
   D_I_175 : FD_732 port map( D => d(175), CK => n49, RESET => n21, Q => Q(175)
                           );
   D_I_176 : FD_731 port map( D => d(176), CK => n50, RESET => n21, Q => Q(176)
                           );
   D_I_177 : FD_730 port map( D => d(177), CK => n50, RESET => n21, Q => Q(177)
                           );
   D_I_178 : FD_729 port map( D => d(178), CK => n50, RESET => n21, Q => Q(178)
                           );
   D_I_179 : FD_728 port map( D => d(179), CK => n50, RESET => n21, Q => Q(179)
                           );
   D_I_180 : FD_727 port map( D => d(180), CK => n50, RESET => n22, Q => Q(180)
                           );
   D_I_181 : FD_726 port map( D => d(181), CK => n50, RESET => n22, Q => Q(181)
                           );
   D_I_182 : FD_725 port map( D => d(182), CK => n50, RESET => n22, Q => Q(182)
                           );
   D_I_183 : FD_724 port map( D => d(183), CK => n50, RESET => n22, Q => Q(183)
                           );
   D_I_184 : FD_723 port map( D => d(184), CK => n50, RESET => n22, Q => Q(184)
                           );
   D_I_185 : FD_722 port map( D => d(185), CK => n50, RESET => n22, Q => Q(185)
                           );
   D_I_186 : FD_721 port map( D => d(186), CK => n50, RESET => n22, Q => Q(186)
                           );
   D_I_187 : FD_720 port map( D => d(187), CK => n51, RESET => n22, Q => Q(187)
                           );
   D_I_188 : FD_719 port map( D => d(188), CK => n51, RESET => n22, Q => Q(188)
                           );
   D_I_189 : FD_718 port map( D => d(189), CK => n51, RESET => n22, Q => Q(189)
                           );
   D_I_190 : FD_717 port map( D => d(190), CK => n51, RESET => n22, Q => Q(190)
                           );
   D_I_191 : FD_716 port map( D => d(191), CK => n51, RESET => n22, Q => Q(191)
                           );
   D_I_192 : FD_715 port map( D => d(192), CK => n51, RESET => n23, Q => Q(192)
                           );
   D_I_193 : FD_714 port map( D => d(193), CK => n51, RESET => n23, Q => Q(193)
                           );
   D_I_194 : FD_713 port map( D => d(194), CK => n51, RESET => n23, Q => Q(194)
                           );
   D_I_195 : FD_712 port map( D => d(195), CK => n51, RESET => n23, Q => Q(195)
                           );
   D_I_196 : FD_711 port map( D => d(196), CK => n51, RESET => n23, Q => Q(196)
                           );
   D_I_197 : FD_710 port map( D => d(197), CK => n51, RESET => n23, Q => Q(197)
                           );
   D_I_198 : FD_709 port map( D => d(198), CK => n52, RESET => n23, Q => Q(198)
                           );
   D_I_199 : FD_708 port map( D => d(199), CK => n52, RESET => n23, Q => Q(199)
                           );
   D_I_200 : FD_707 port map( D => d(200), CK => n52, RESET => n23, Q => Q(200)
                           );
   D_I_201 : FD_706 port map( D => d(201), CK => n52, RESET => n23, Q => Q(201)
                           );
   D_I_202 : FD_705 port map( D => d(202), CK => n52, RESET => n23, Q => Q(202)
                           );
   D_I_203 : FD_704 port map( D => d(203), CK => n52, RESET => n23, Q => Q(203)
                           );
   D_I_204 : FD_703 port map( D => d(204), CK => n52, RESET => n24, Q => Q(204)
                           );
   D_I_205 : FD_702 port map( D => d(205), CK => n52, RESET => n24, Q => Q(205)
                           );
   D_I_206 : FD_701 port map( D => d(206), CK => n52, RESET => n24, Q => Q(206)
                           );
   D_I_207 : FD_700 port map( D => d(207), CK => n52, RESET => n24, Q => Q(207)
                           );
   D_I_208 : FD_699 port map( D => d(208), CK => n52, RESET => n24, Q => Q(208)
                           );
   D_I_209 : FD_698 port map( D => d(209), CK => n53, RESET => n24, Q => Q(209)
                           );
   D_I_210 : FD_697 port map( D => d(210), CK => n53, RESET => n24, Q => Q(210)
                           );
   D_I_211 : FD_696 port map( D => d(211), CK => n53, RESET => n24, Q => Q(211)
                           );
   D_I_212 : FD_695 port map( D => d(212), CK => n53, RESET => n24, Q => Q(212)
                           );
   D_I_213 : FD_694 port map( D => d(213), CK => n53, RESET => n24, Q => Q(213)
                           );
   D_I_214 : FD_693 port map( D => d(214), CK => n53, RESET => n24, Q => Q(214)
                           );
   D_I_215 : FD_692 port map( D => d(215), CK => n53, RESET => n24, Q => Q(215)
                           );
   D_I_216 : FD_691 port map( D => d(216), CK => n53, RESET => n25, Q => Q(216)
                           );
   D_I_217 : FD_690 port map( D => d(217), CK => n53, RESET => n25, Q => Q(217)
                           );
   D_I_218 : FD_689 port map( D => d(218), CK => n53, RESET => n25, Q => Q(218)
                           );
   D_I_219 : FD_688 port map( D => d(219), CK => n53, RESET => n25, Q => Q(219)
                           );
   D_I_220 : FD_687 port map( D => d(220), CK => n54, RESET => n25, Q => Q(220)
                           );
   D_I_221 : FD_686 port map( D => d(221), CK => n54, RESET => n25, Q => Q(221)
                           );
   D_I_222 : FD_685 port map( D => d(222), CK => n54, RESET => n25, Q => Q(222)
                           );
   D_I_223 : FD_684 port map( D => d(223), CK => n54, RESET => n25, Q => Q(223)
                           );
   D_I_224 : FD_683 port map( D => d(224), CK => n54, RESET => n25, Q => Q(224)
                           );
   D_I_225 : FD_682 port map( D => d(225), CK => n54, RESET => n25, Q => Q(225)
                           );
   D_I_226 : FD_681 port map( D => d(226), CK => n54, RESET => n25, Q => Q(226)
                           );
   D_I_227 : FD_680 port map( D => d(227), CK => n54, RESET => n25, Q => Q(227)
                           );
   D_I_228 : FD_679 port map( D => d(228), CK => n54, RESET => n26, Q => Q(228)
                           );
   D_I_229 : FD_678 port map( D => d(229), CK => n54, RESET => n26, Q => Q(229)
                           );
   D_I_230 : FD_677 port map( D => d(230), CK => n54, RESET => n26, Q => Q(230)
                           );
   D_I_231 : FD_676 port map( D => d(231), CK => n55, RESET => n26, Q => Q(231)
                           );
   D_I_232 : FD_675 port map( D => d(232), CK => n55, RESET => n26, Q => Q(232)
                           );
   D_I_233 : FD_674 port map( D => d(233), CK => n55, RESET => n26, Q => Q(233)
                           );
   D_I_234 : FD_673 port map( D => d(234), CK => n55, RESET => n26, Q => Q(234)
                           );
   D_I_235 : FD_672 port map( D => d(235), CK => n55, RESET => n26, Q => Q(235)
                           );
   D_I_236 : FD_671 port map( D => d(236), CK => n55, RESET => n26, Q => Q(236)
                           );
   D_I_237 : FD_670 port map( D => d(237), CK => n55, RESET => n26, Q => Q(237)
                           );
   D_I_238 : FD_669 port map( D => d(238), CK => n55, RESET => n26, Q => Q(238)
                           );
   D_I_239 : FD_668 port map( D => d(239), CK => n55, RESET => n26, Q => Q(239)
                           );
   D_I_240 : FD_667 port map( D => d(240), CK => n55, RESET => n27, Q => Q(240)
                           );
   D_I_241 : FD_666 port map( D => d(241), CK => n55, RESET => n27, Q => Q(241)
                           );
   D_I_242 : FD_665 port map( D => d(242), CK => n56, RESET => n27, Q => Q(242)
                           );
   D_I_243 : FD_664 port map( D => d(243), CK => n56, RESET => n27, Q => Q(243)
                           );
   D_I_244 : FD_663 port map( D => d(244), CK => n56, RESET => n27, Q => Q(244)
                           );
   D_I_245 : FD_662 port map( D => d(245), CK => n56, RESET => n27, Q => Q(245)
                           );
   D_I_246 : FD_661 port map( D => d(246), CK => n56, RESET => n27, Q => Q(246)
                           );
   D_I_247 : FD_660 port map( D => d(247), CK => n56, RESET => n27, Q => Q(247)
                           );
   D_I_248 : FD_659 port map( D => d(248), CK => n56, RESET => n27, Q => Q(248)
                           );
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_2 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_2;

architecture SYN_struc of reg_nbit_n249_2 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_378
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_379
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_380
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_381
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_382
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_383
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_384
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_385
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_386
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_387
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_388
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_389
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_390
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_391
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_392
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_393
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_394
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_395
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_396
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_397
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_398
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_399
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_400
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_401
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_402
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_403
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_404
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_405
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_406
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_407
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_408
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_409
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_410
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_411
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_412
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_413
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_414
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_415
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_416
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_417
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_418
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_419
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_420
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_421
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_422
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_423
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_424
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_425
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_426
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_427
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_428
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_429
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_430
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_431
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_432
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_433
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_434
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_435
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_436
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_437
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_438
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_439
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_440
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_441
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_442
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_443
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_444
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_445
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_446
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_447
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_448
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_449
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_450
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_451
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_452
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_453
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_454
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_455
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_456
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_457
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_458
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_459
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_460
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_461
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_462
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_463
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_464
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_465
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_466
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_467
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_468
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_469
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_470
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_471
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_472
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_473
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_474
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_475
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_476
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_477
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_478
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_479
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_480
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_481
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_482
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_483
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_484
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_485
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_486
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_487
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_488
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_489
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_490
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_491
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_492
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_493
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_494
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_495
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_496
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_497
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_498
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_499
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_500
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_501
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_502
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_503
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_504
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_505
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_506
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_507
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_508
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_509
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_510
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_511
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_512
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_513
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_514
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_515
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_516
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_517
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_518
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_519
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_520
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_521
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_522
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_523
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_524
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_525
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_526
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_527
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_528
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_529
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_530
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_531
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_532
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_533
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_534
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_535
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_536
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_537
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_538
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_539
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_540
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_541
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_542
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_543
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_544
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_545
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_546
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_547
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_548
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_549
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_550
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_551
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_552
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_553
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_554
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_555
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_556
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_557
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_558
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_559
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_560
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_561
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_562
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_563
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_564
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_565
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_566
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_567
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_568
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_569
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_570
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_571
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_572
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_573
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_574
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_575
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_576
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_577
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_578
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_579
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_580
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_581
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_582
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_583
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_584
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_585
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_586
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_587
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_588
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_589
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_590
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_591
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_592
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_593
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_594
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_595
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_596
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_597
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_598
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_599
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_600
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_601
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_602
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_603
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_604
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_605
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_606
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_607
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_608
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_609
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_610
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_611
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_612
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_613
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_614
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_615
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_616
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_617
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_618
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_619
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_620
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_621
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_622
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_623
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_624
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_625
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_626
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_626 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_625 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_624 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_623 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_622 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_621 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_620 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_619 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_618 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_617 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_616 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_615 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_614 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_613 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_612 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_611 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_610 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_609 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_608 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_607 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_606 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_605 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_604 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_603 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_602 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_601 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_600 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_599 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_598 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_597 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_596 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_595 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_594 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_593 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_592 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_591 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_590 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_589 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_588 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_587 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_586 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_585 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_584 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_583 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_582 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_581 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_580 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_579 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_578 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_577 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_576 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_575 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_574 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_573 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_572 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_571 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_570 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_569 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_568 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_567 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_566 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_565 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_564 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_563 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_562 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_561 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_560 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_559 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_558 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_557 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_556 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_555 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_554 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_553 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_552 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_551 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_550 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_549 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_548 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_547 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_546 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_545 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_544 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_543 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_542 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_541 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_540 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_539 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_538 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_537 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_536 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_535 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_534 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_533 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_532 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_531 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_530 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_529 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_528 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_527 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_526 port map( D => d(100), CK => n43, RESET => n15, Q => Q(100)
                           );
   D_I_101 : FD_525 port map( D => d(101), CK => n43, RESET => n15, Q => Q(101)
                           );
   D_I_102 : FD_524 port map( D => d(102), CK => n43, RESET => n15, Q => Q(102)
                           );
   D_I_103 : FD_523 port map( D => d(103), CK => n43, RESET => n15, Q => Q(103)
                           );
   D_I_104 : FD_522 port map( D => d(104), CK => n43, RESET => n15, Q => Q(104)
                           );
   D_I_105 : FD_521 port map( D => d(105), CK => n43, RESET => n15, Q => Q(105)
                           );
   D_I_106 : FD_520 port map( D => d(106), CK => n43, RESET => n15, Q => Q(106)
                           );
   D_I_107 : FD_519 port map( D => d(107), CK => n43, RESET => n15, Q => Q(107)
                           );
   D_I_108 : FD_518 port map( D => d(108), CK => n43, RESET => n16, Q => Q(108)
                           );
   D_I_109 : FD_517 port map( D => d(109), CK => n43, RESET => n16, Q => Q(109)
                           );
   D_I_110 : FD_516 port map( D => d(110), CK => n44, RESET => n16, Q => Q(110)
                           );
   D_I_111 : FD_515 port map( D => d(111), CK => n44, RESET => n16, Q => Q(111)
                           );
   D_I_112 : FD_514 port map( D => d(112), CK => n44, RESET => n16, Q => Q(112)
                           );
   D_I_113 : FD_513 port map( D => d(113), CK => n44, RESET => n16, Q => Q(113)
                           );
   D_I_114 : FD_512 port map( D => d(114), CK => n44, RESET => n16, Q => Q(114)
                           );
   D_I_115 : FD_511 port map( D => d(115), CK => n44, RESET => n16, Q => Q(115)
                           );
   D_I_116 : FD_510 port map( D => d(116), CK => n44, RESET => n16, Q => Q(116)
                           );
   D_I_117 : FD_509 port map( D => d(117), CK => n44, RESET => n16, Q => Q(117)
                           );
   D_I_118 : FD_508 port map( D => d(118), CK => n44, RESET => n16, Q => Q(118)
                           );
   D_I_119 : FD_507 port map( D => d(119), CK => n44, RESET => n16, Q => Q(119)
                           );
   D_I_120 : FD_506 port map( D => d(120), CK => n44, RESET => n17, Q => Q(120)
                           );
   D_I_121 : FD_505 port map( D => d(121), CK => n45, RESET => n17, Q => Q(121)
                           );
   D_I_122 : FD_504 port map( D => d(122), CK => n45, RESET => n17, Q => Q(122)
                           );
   D_I_123 : FD_503 port map( D => d(123), CK => n45, RESET => n17, Q => Q(123)
                           );
   D_I_124 : FD_502 port map( D => d(124), CK => n45, RESET => n17, Q => Q(124)
                           );
   D_I_125 : FD_501 port map( D => d(125), CK => n45, RESET => n17, Q => Q(125)
                           );
   D_I_126 : FD_500 port map( D => d(126), CK => n45, RESET => n17, Q => Q(126)
                           );
   D_I_127 : FD_499 port map( D => d(127), CK => n45, RESET => n17, Q => Q(127)
                           );
   D_I_128 : FD_498 port map( D => d(128), CK => n45, RESET => n17, Q => Q(128)
                           );
   D_I_129 : FD_497 port map( D => d(129), CK => n45, RESET => n17, Q => Q(129)
                           );
   D_I_130 : FD_496 port map( D => d(130), CK => n45, RESET => n17, Q => Q(130)
                           );
   D_I_131 : FD_495 port map( D => d(131), CK => n45, RESET => n17, Q => Q(131)
                           );
   D_I_132 : FD_494 port map( D => d(132), CK => n46, RESET => n18, Q => Q(132)
                           );
   D_I_133 : FD_493 port map( D => d(133), CK => n46, RESET => n18, Q => Q(133)
                           );
   D_I_134 : FD_492 port map( D => d(134), CK => n46, RESET => n18, Q => Q(134)
                           );
   D_I_135 : FD_491 port map( D => d(135), CK => n46, RESET => n18, Q => Q(135)
                           );
   D_I_136 : FD_490 port map( D => d(136), CK => n46, RESET => n18, Q => Q(136)
                           );
   D_I_137 : FD_489 port map( D => d(137), CK => n46, RESET => n18, Q => Q(137)
                           );
   D_I_138 : FD_488 port map( D => d(138), CK => n46, RESET => n18, Q => Q(138)
                           );
   D_I_139 : FD_487 port map( D => d(139), CK => n46, RESET => n18, Q => Q(139)
                           );
   D_I_140 : FD_486 port map( D => d(140), CK => n46, RESET => n18, Q => Q(140)
                           );
   D_I_141 : FD_485 port map( D => d(141), CK => n46, RESET => n18, Q => Q(141)
                           );
   D_I_142 : FD_484 port map( D => d(142), CK => n46, RESET => n18, Q => Q(142)
                           );
   D_I_143 : FD_483 port map( D => d(143), CK => n47, RESET => n18, Q => Q(143)
                           );
   D_I_144 : FD_482 port map( D => d(144), CK => n47, RESET => n19, Q => Q(144)
                           );
   D_I_145 : FD_481 port map( D => d(145), CK => n47, RESET => n19, Q => Q(145)
                           );
   D_I_146 : FD_480 port map( D => d(146), CK => n47, RESET => n19, Q => Q(146)
                           );
   D_I_147 : FD_479 port map( D => d(147), CK => n47, RESET => n19, Q => Q(147)
                           );
   D_I_148 : FD_478 port map( D => d(148), CK => n47, RESET => n19, Q => Q(148)
                           );
   D_I_149 : FD_477 port map( D => d(149), CK => n47, RESET => n19, Q => Q(149)
                           );
   D_I_150 : FD_476 port map( D => d(150), CK => n47, RESET => n19, Q => Q(150)
                           );
   D_I_151 : FD_475 port map( D => d(151), CK => n47, RESET => n19, Q => Q(151)
                           );
   D_I_152 : FD_474 port map( D => d(152), CK => n47, RESET => n19, Q => Q(152)
                           );
   D_I_153 : FD_473 port map( D => d(153), CK => n47, RESET => n19, Q => Q(153)
                           );
   D_I_154 : FD_472 port map( D => d(154), CK => n48, RESET => n19, Q => Q(154)
                           );
   D_I_155 : FD_471 port map( D => d(155), CK => n48, RESET => n19, Q => Q(155)
                           );
   D_I_156 : FD_470 port map( D => d(156), CK => n48, RESET => n20, Q => Q(156)
                           );
   D_I_157 : FD_469 port map( D => d(157), CK => n48, RESET => n20, Q => Q(157)
                           );
   D_I_158 : FD_468 port map( D => d(158), CK => n48, RESET => n20, Q => Q(158)
                           );
   D_I_159 : FD_467 port map( D => d(159), CK => n48, RESET => n20, Q => Q(159)
                           );
   D_I_160 : FD_466 port map( D => d(160), CK => n48, RESET => n20, Q => Q(160)
                           );
   D_I_161 : FD_465 port map( D => d(161), CK => n48, RESET => n20, Q => Q(161)
                           );
   D_I_162 : FD_464 port map( D => d(162), CK => n48, RESET => n20, Q => Q(162)
                           );
   D_I_163 : FD_463 port map( D => d(163), CK => n48, RESET => n20, Q => Q(163)
                           );
   D_I_164 : FD_462 port map( D => d(164), CK => n48, RESET => n20, Q => Q(164)
                           );
   D_I_165 : FD_461 port map( D => d(165), CK => n49, RESET => n20, Q => Q(165)
                           );
   D_I_166 : FD_460 port map( D => d(166), CK => n49, RESET => n20, Q => Q(166)
                           );
   D_I_167 : FD_459 port map( D => d(167), CK => n49, RESET => n20, Q => Q(167)
                           );
   D_I_168 : FD_458 port map( D => d(168), CK => n49, RESET => n21, Q => Q(168)
                           );
   D_I_169 : FD_457 port map( D => d(169), CK => n49, RESET => n21, Q => Q(169)
                           );
   D_I_170 : FD_456 port map( D => d(170), CK => n49, RESET => n21, Q => Q(170)
                           );
   D_I_171 : FD_455 port map( D => d(171), CK => n49, RESET => n21, Q => Q(171)
                           );
   D_I_172 : FD_454 port map( D => d(172), CK => n49, RESET => n21, Q => Q(172)
                           );
   D_I_173 : FD_453 port map( D => d(173), CK => n49, RESET => n21, Q => Q(173)
                           );
   D_I_174 : FD_452 port map( D => d(174), CK => n49, RESET => n21, Q => Q(174)
                           );
   D_I_175 : FD_451 port map( D => d(175), CK => n49, RESET => n21, Q => Q(175)
                           );
   D_I_176 : FD_450 port map( D => d(176), CK => n50, RESET => n21, Q => Q(176)
                           );
   D_I_177 : FD_449 port map( D => d(177), CK => n50, RESET => n21, Q => Q(177)
                           );
   D_I_178 : FD_448 port map( D => d(178), CK => n50, RESET => n21, Q => Q(178)
                           );
   D_I_179 : FD_447 port map( D => d(179), CK => n50, RESET => n21, Q => Q(179)
                           );
   D_I_180 : FD_446 port map( D => d(180), CK => n50, RESET => n22, Q => Q(180)
                           );
   D_I_181 : FD_445 port map( D => d(181), CK => n50, RESET => n22, Q => Q(181)
                           );
   D_I_182 : FD_444 port map( D => d(182), CK => n50, RESET => n22, Q => Q(182)
                           );
   D_I_183 : FD_443 port map( D => d(183), CK => n50, RESET => n22, Q => Q(183)
                           );
   D_I_184 : FD_442 port map( D => d(184), CK => n50, RESET => n22, Q => Q(184)
                           );
   D_I_185 : FD_441 port map( D => d(185), CK => n50, RESET => n22, Q => Q(185)
                           );
   D_I_186 : FD_440 port map( D => d(186), CK => n50, RESET => n22, Q => Q(186)
                           );
   D_I_187 : FD_439 port map( D => d(187), CK => n51, RESET => n22, Q => Q(187)
                           );
   D_I_188 : FD_438 port map( D => d(188), CK => n51, RESET => n22, Q => Q(188)
                           );
   D_I_189 : FD_437 port map( D => d(189), CK => n51, RESET => n22, Q => Q(189)
                           );
   D_I_190 : FD_436 port map( D => d(190), CK => n51, RESET => n22, Q => Q(190)
                           );
   D_I_191 : FD_435 port map( D => d(191), CK => n51, RESET => n22, Q => Q(191)
                           );
   D_I_192 : FD_434 port map( D => d(192), CK => n51, RESET => n23, Q => Q(192)
                           );
   D_I_193 : FD_433 port map( D => d(193), CK => n51, RESET => n23, Q => Q(193)
                           );
   D_I_194 : FD_432 port map( D => d(194), CK => n51, RESET => n23, Q => Q(194)
                           );
   D_I_195 : FD_431 port map( D => d(195), CK => n51, RESET => n23, Q => Q(195)
                           );
   D_I_196 : FD_430 port map( D => d(196), CK => n51, RESET => n23, Q => Q(196)
                           );
   D_I_197 : FD_429 port map( D => d(197), CK => n51, RESET => n23, Q => Q(197)
                           );
   D_I_198 : FD_428 port map( D => d(198), CK => n52, RESET => n23, Q => Q(198)
                           );
   D_I_199 : FD_427 port map( D => d(199), CK => n52, RESET => n23, Q => Q(199)
                           );
   D_I_200 : FD_426 port map( D => d(200), CK => n52, RESET => n23, Q => Q(200)
                           );
   D_I_201 : FD_425 port map( D => d(201), CK => n52, RESET => n23, Q => Q(201)
                           );
   D_I_202 : FD_424 port map( D => d(202), CK => n52, RESET => n23, Q => Q(202)
                           );
   D_I_203 : FD_423 port map( D => d(203), CK => n52, RESET => n23, Q => Q(203)
                           );
   D_I_204 : FD_422 port map( D => d(204), CK => n52, RESET => n24, Q => Q(204)
                           );
   D_I_205 : FD_421 port map( D => d(205), CK => n52, RESET => n24, Q => Q(205)
                           );
   D_I_206 : FD_420 port map( D => d(206), CK => n52, RESET => n24, Q => Q(206)
                           );
   D_I_207 : FD_419 port map( D => d(207), CK => n52, RESET => n24, Q => Q(207)
                           );
   D_I_208 : FD_418 port map( D => d(208), CK => n52, RESET => n24, Q => Q(208)
                           );
   D_I_209 : FD_417 port map( D => d(209), CK => n53, RESET => n24, Q => Q(209)
                           );
   D_I_210 : FD_416 port map( D => d(210), CK => n53, RESET => n24, Q => Q(210)
                           );
   D_I_211 : FD_415 port map( D => d(211), CK => n53, RESET => n24, Q => Q(211)
                           );
   D_I_212 : FD_414 port map( D => d(212), CK => n53, RESET => n24, Q => Q(212)
                           );
   D_I_213 : FD_413 port map( D => d(213), CK => n53, RESET => n24, Q => Q(213)
                           );
   D_I_214 : FD_412 port map( D => d(214), CK => n53, RESET => n24, Q => Q(214)
                           );
   D_I_215 : FD_411 port map( D => d(215), CK => n53, RESET => n24, Q => Q(215)
                           );
   D_I_216 : FD_410 port map( D => d(216), CK => n53, RESET => n25, Q => Q(216)
                           );
   D_I_217 : FD_409 port map( D => d(217), CK => n53, RESET => n25, Q => Q(217)
                           );
   D_I_218 : FD_408 port map( D => d(218), CK => n53, RESET => n25, Q => Q(218)
                           );
   D_I_219 : FD_407 port map( D => d(219), CK => n53, RESET => n25, Q => Q(219)
                           );
   D_I_220 : FD_406 port map( D => d(220), CK => n54, RESET => n25, Q => Q(220)
                           );
   D_I_221 : FD_405 port map( D => d(221), CK => n54, RESET => n25, Q => Q(221)
                           );
   D_I_222 : FD_404 port map( D => d(222), CK => n54, RESET => n25, Q => Q(222)
                           );
   D_I_223 : FD_403 port map( D => d(223), CK => n54, RESET => n25, Q => Q(223)
                           );
   D_I_224 : FD_402 port map( D => d(224), CK => n54, RESET => n25, Q => Q(224)
                           );
   D_I_225 : FD_401 port map( D => d(225), CK => n54, RESET => n25, Q => Q(225)
                           );
   D_I_226 : FD_400 port map( D => d(226), CK => n54, RESET => n25, Q => Q(226)
                           );
   D_I_227 : FD_399 port map( D => d(227), CK => n54, RESET => n25, Q => Q(227)
                           );
   D_I_228 : FD_398 port map( D => d(228), CK => n54, RESET => n26, Q => Q(228)
                           );
   D_I_229 : FD_397 port map( D => d(229), CK => n54, RESET => n26, Q => Q(229)
                           );
   D_I_230 : FD_396 port map( D => d(230), CK => n54, RESET => n26, Q => Q(230)
                           );
   D_I_231 : FD_395 port map( D => d(231), CK => n55, RESET => n26, Q => Q(231)
                           );
   D_I_232 : FD_394 port map( D => d(232), CK => n55, RESET => n26, Q => Q(232)
                           );
   D_I_233 : FD_393 port map( D => d(233), CK => n55, RESET => n26, Q => Q(233)
                           );
   D_I_234 : FD_392 port map( D => d(234), CK => n55, RESET => n26, Q => Q(234)
                           );
   D_I_235 : FD_391 port map( D => d(235), CK => n55, RESET => n26, Q => Q(235)
                           );
   D_I_236 : FD_390 port map( D => d(236), CK => n55, RESET => n26, Q => Q(236)
                           );
   D_I_237 : FD_389 port map( D => d(237), CK => n55, RESET => n26, Q => Q(237)
                           );
   D_I_238 : FD_388 port map( D => d(238), CK => n55, RESET => n26, Q => Q(238)
                           );
   D_I_239 : FD_387 port map( D => d(239), CK => n55, RESET => n26, Q => Q(239)
                           );
   D_I_240 : FD_386 port map( D => d(240), CK => n55, RESET => n27, Q => Q(240)
                           );
   D_I_241 : FD_385 port map( D => d(241), CK => n55, RESET => n27, Q => Q(241)
                           );
   D_I_242 : FD_384 port map( D => d(242), CK => n56, RESET => n27, Q => Q(242)
                           );
   D_I_243 : FD_383 port map( D => d(243), CK => n56, RESET => n27, Q => Q(243)
                           );
   D_I_244 : FD_382 port map( D => d(244), CK => n56, RESET => n27, Q => Q(244)
                           );
   D_I_245 : FD_381 port map( D => d(245), CK => n56, RESET => n27, Q => Q(245)
                           );
   D_I_246 : FD_380 port map( D => d(246), CK => n56, RESET => n27, Q => Q(246)
                           );
   D_I_247 : FD_379 port map( D => d(247), CK => n56, RESET => n27, Q => Q(247)
                           );
   D_I_248 : FD_378 port map( D => d(248), CK => n56, RESET => n27, Q => Q(248)
                           );
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_1;

architecture SYN_struc of reg_nbit_n249_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_97
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_98
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_99
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_100
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_101
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_102
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_103
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_104
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_105
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_106
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_107
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_108
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_109
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_110
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_111
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_112
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_113
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_114
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_115
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_116
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_117
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_118
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_119
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_120
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_121
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_122
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_123
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_124
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_125
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_126
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_127
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_128
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_129
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_130
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_131
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_132
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_133
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_134
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_135
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_136
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_137
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_138
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_139
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_140
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_141
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_142
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_143
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_144
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_145
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_146
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_147
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_148
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_149
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_150
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_151
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_152
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_153
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_154
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_155
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_156
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_157
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_158
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_159
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_160
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_161
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_162
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_163
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_164
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_165
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_166
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_167
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_168
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_169
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_170
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_171
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_172
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_173
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_174
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_175
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_176
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_177
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_178
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_179
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_180
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_181
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_182
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_183
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_184
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_185
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_186
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_187
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_188
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_189
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_190
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_191
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_192
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_193
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_194
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_195
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_196
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_197
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_198
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_199
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_200
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_201
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_202
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_203
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_204
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_205
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_206
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_207
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_208
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_209
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_210
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_211
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_212
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_213
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_214
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_215
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_216
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_217
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_218
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_219
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_220
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_221
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_222
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_223
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_224
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_225
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_226
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_227
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_228
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_229
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_230
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_231
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_232
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_233
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_234
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_235
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_236
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_237
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_238
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_239
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_240
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_241
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_242
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_243
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_244
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_245
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_246
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_247
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_248
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_249
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_250
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_251
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_252
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_253
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_254
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_255
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_256
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_257
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_258
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_259
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_260
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_261
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_262
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_263
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_264
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_265
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_266
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_267
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_268
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_269
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_270
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_271
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_272
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_273
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_274
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_275
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_276
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_277
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_278
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_279
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_280
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_281
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_282
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_283
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_284
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_285
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_286
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_287
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_288
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_289
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_290
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_291
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_292
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_293
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_294
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_295
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_296
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_297
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_298
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_299
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_300
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_301
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_302
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_303
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_304
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_305
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_306
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_307
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_308
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_309
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_310
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_311
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_312
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_313
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_314
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_315
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_316
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_317
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_318
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_319
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_320
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_321
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_322
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_323
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_324
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_325
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_326
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_327
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_328
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_329
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_330
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_331
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_332
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_333
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_334
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_335
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_336
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_337
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_338
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_339
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_340
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_341
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_342
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_343
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_344
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_345
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_345 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_344 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_343 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_342 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_341 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_340 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_339 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_338 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_337 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_336 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_335 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_334 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_333 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_332 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_331 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_330 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_329 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_328 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_327 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_326 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_325 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_324 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_323 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_322 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_321 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_320 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_319 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_318 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_317 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_316 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_315 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_314 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_313 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_312 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_311 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_310 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_309 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_308 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_307 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_306 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_305 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_304 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_303 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_302 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_301 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_300 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_299 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_298 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_297 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_296 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_295 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_294 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_293 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_292 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_291 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_290 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_289 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_288 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_287 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_286 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_285 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_284 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_283 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_282 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_281 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_280 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_279 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_278 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_277 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_276 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_275 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_274 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_273 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_272 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_271 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_270 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_269 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_268 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_267 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_266 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_265 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_264 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_263 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_262 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_261 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_260 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_259 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_258 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_257 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_256 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_255 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_254 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_253 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_252 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_251 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_250 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_249 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_248 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_247 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_246 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_245 port map( D => d(100), CK => n43, RESET => n15, Q => Q(100)
                           );
   D_I_101 : FD_244 port map( D => d(101), CK => n43, RESET => n15, Q => Q(101)
                           );
   D_I_102 : FD_243 port map( D => d(102), CK => n43, RESET => n15, Q => Q(102)
                           );
   D_I_103 : FD_242 port map( D => d(103), CK => n43, RESET => n15, Q => Q(103)
                           );
   D_I_104 : FD_241 port map( D => d(104), CK => n43, RESET => n15, Q => Q(104)
                           );
   D_I_105 : FD_240 port map( D => d(105), CK => n43, RESET => n15, Q => Q(105)
                           );
   D_I_106 : FD_239 port map( D => d(106), CK => n43, RESET => n15, Q => Q(106)
                           );
   D_I_107 : FD_238 port map( D => d(107), CK => n43, RESET => n15, Q => Q(107)
                           );
   D_I_108 : FD_237 port map( D => d(108), CK => n43, RESET => n16, Q => Q(108)
                           );
   D_I_109 : FD_236 port map( D => d(109), CK => n43, RESET => n16, Q => Q(109)
                           );
   D_I_110 : FD_235 port map( D => d(110), CK => n44, RESET => n16, Q => Q(110)
                           );
   D_I_111 : FD_234 port map( D => d(111), CK => n44, RESET => n16, Q => Q(111)
                           );
   D_I_112 : FD_233 port map( D => d(112), CK => n44, RESET => n16, Q => Q(112)
                           );
   D_I_113 : FD_232 port map( D => d(113), CK => n44, RESET => n16, Q => Q(113)
                           );
   D_I_114 : FD_231 port map( D => d(114), CK => n44, RESET => n16, Q => Q(114)
                           );
   D_I_115 : FD_230 port map( D => d(115), CK => n44, RESET => n16, Q => Q(115)
                           );
   D_I_116 : FD_229 port map( D => d(116), CK => n44, RESET => n16, Q => Q(116)
                           );
   D_I_117 : FD_228 port map( D => d(117), CK => n44, RESET => n16, Q => Q(117)
                           );
   D_I_118 : FD_227 port map( D => d(118), CK => n44, RESET => n16, Q => Q(118)
                           );
   D_I_119 : FD_226 port map( D => d(119), CK => n44, RESET => n16, Q => Q(119)
                           );
   D_I_120 : FD_225 port map( D => d(120), CK => n44, RESET => n17, Q => Q(120)
                           );
   D_I_121 : FD_224 port map( D => d(121), CK => n45, RESET => n17, Q => Q(121)
                           );
   D_I_122 : FD_223 port map( D => d(122), CK => n45, RESET => n17, Q => Q(122)
                           );
   D_I_123 : FD_222 port map( D => d(123), CK => n45, RESET => n17, Q => Q(123)
                           );
   D_I_124 : FD_221 port map( D => d(124), CK => n45, RESET => n17, Q => Q(124)
                           );
   D_I_125 : FD_220 port map( D => d(125), CK => n45, RESET => n17, Q => Q(125)
                           );
   D_I_126 : FD_219 port map( D => d(126), CK => n45, RESET => n17, Q => Q(126)
                           );
   D_I_127 : FD_218 port map( D => d(127), CK => n45, RESET => n17, Q => Q(127)
                           );
   D_I_128 : FD_217 port map( D => d(128), CK => n45, RESET => n17, Q => Q(128)
                           );
   D_I_129 : FD_216 port map( D => d(129), CK => n45, RESET => n17, Q => Q(129)
                           );
   D_I_130 : FD_215 port map( D => d(130), CK => n45, RESET => n17, Q => Q(130)
                           );
   D_I_131 : FD_214 port map( D => d(131), CK => n45, RESET => n17, Q => Q(131)
                           );
   D_I_132 : FD_213 port map( D => d(132), CK => n46, RESET => n18, Q => Q(132)
                           );
   D_I_133 : FD_212 port map( D => d(133), CK => n46, RESET => n18, Q => Q(133)
                           );
   D_I_134 : FD_211 port map( D => d(134), CK => n46, RESET => n18, Q => Q(134)
                           );
   D_I_135 : FD_210 port map( D => d(135), CK => n46, RESET => n18, Q => Q(135)
                           );
   D_I_136 : FD_209 port map( D => d(136), CK => n46, RESET => n18, Q => Q(136)
                           );
   D_I_137 : FD_208 port map( D => d(137), CK => n46, RESET => n18, Q => Q(137)
                           );
   D_I_138 : FD_207 port map( D => d(138), CK => n46, RESET => n18, Q => Q(138)
                           );
   D_I_139 : FD_206 port map( D => d(139), CK => n46, RESET => n18, Q => Q(139)
                           );
   D_I_140 : FD_205 port map( D => d(140), CK => n46, RESET => n18, Q => Q(140)
                           );
   D_I_141 : FD_204 port map( D => d(141), CK => n46, RESET => n18, Q => Q(141)
                           );
   D_I_142 : FD_203 port map( D => d(142), CK => n46, RESET => n18, Q => Q(142)
                           );
   D_I_143 : FD_202 port map( D => d(143), CK => n47, RESET => n18, Q => Q(143)
                           );
   D_I_144 : FD_201 port map( D => d(144), CK => n47, RESET => n19, Q => Q(144)
                           );
   D_I_145 : FD_200 port map( D => d(145), CK => n47, RESET => n19, Q => Q(145)
                           );
   D_I_146 : FD_199 port map( D => d(146), CK => n47, RESET => n19, Q => Q(146)
                           );
   D_I_147 : FD_198 port map( D => d(147), CK => n47, RESET => n19, Q => Q(147)
                           );
   D_I_148 : FD_197 port map( D => d(148), CK => n47, RESET => n19, Q => Q(148)
                           );
   D_I_149 : FD_196 port map( D => d(149), CK => n47, RESET => n19, Q => Q(149)
                           );
   D_I_150 : FD_195 port map( D => d(150), CK => n47, RESET => n19, Q => Q(150)
                           );
   D_I_151 : FD_194 port map( D => d(151), CK => n47, RESET => n19, Q => Q(151)
                           );
   D_I_152 : FD_193 port map( D => d(152), CK => n47, RESET => n19, Q => Q(152)
                           );
   D_I_153 : FD_192 port map( D => d(153), CK => n47, RESET => n19, Q => Q(153)
                           );
   D_I_154 : FD_191 port map( D => d(154), CK => n48, RESET => n19, Q => Q(154)
                           );
   D_I_155 : FD_190 port map( D => d(155), CK => n48, RESET => n19, Q => Q(155)
                           );
   D_I_156 : FD_189 port map( D => d(156), CK => n48, RESET => n20, Q => Q(156)
                           );
   D_I_157 : FD_188 port map( D => d(157), CK => n48, RESET => n20, Q => Q(157)
                           );
   D_I_158 : FD_187 port map( D => d(158), CK => n48, RESET => n20, Q => Q(158)
                           );
   D_I_159 : FD_186 port map( D => d(159), CK => n48, RESET => n20, Q => Q(159)
                           );
   D_I_160 : FD_185 port map( D => d(160), CK => n48, RESET => n20, Q => Q(160)
                           );
   D_I_161 : FD_184 port map( D => d(161), CK => n48, RESET => n20, Q => Q(161)
                           );
   D_I_162 : FD_183 port map( D => d(162), CK => n48, RESET => n20, Q => Q(162)
                           );
   D_I_163 : FD_182 port map( D => d(163), CK => n48, RESET => n20, Q => Q(163)
                           );
   D_I_164 : FD_181 port map( D => d(164), CK => n48, RESET => n20, Q => Q(164)
                           );
   D_I_165 : FD_180 port map( D => d(165), CK => n49, RESET => n20, Q => Q(165)
                           );
   D_I_166 : FD_179 port map( D => d(166), CK => n49, RESET => n20, Q => Q(166)
                           );
   D_I_167 : FD_178 port map( D => d(167), CK => n49, RESET => n20, Q => Q(167)
                           );
   D_I_168 : FD_177 port map( D => d(168), CK => n49, RESET => n21, Q => Q(168)
                           );
   D_I_169 : FD_176 port map( D => d(169), CK => n49, RESET => n21, Q => Q(169)
                           );
   D_I_170 : FD_175 port map( D => d(170), CK => n49, RESET => n21, Q => Q(170)
                           );
   D_I_171 : FD_174 port map( D => d(171), CK => n49, RESET => n21, Q => Q(171)
                           );
   D_I_172 : FD_173 port map( D => d(172), CK => n49, RESET => n21, Q => Q(172)
                           );
   D_I_173 : FD_172 port map( D => d(173), CK => n49, RESET => n21, Q => Q(173)
                           );
   D_I_174 : FD_171 port map( D => d(174), CK => n49, RESET => n21, Q => Q(174)
                           );
   D_I_175 : FD_170 port map( D => d(175), CK => n49, RESET => n21, Q => Q(175)
                           );
   D_I_176 : FD_169 port map( D => d(176), CK => n50, RESET => n21, Q => Q(176)
                           );
   D_I_177 : FD_168 port map( D => d(177), CK => n50, RESET => n21, Q => Q(177)
                           );
   D_I_178 : FD_167 port map( D => d(178), CK => n50, RESET => n21, Q => Q(178)
                           );
   D_I_179 : FD_166 port map( D => d(179), CK => n50, RESET => n21, Q => Q(179)
                           );
   D_I_180 : FD_165 port map( D => d(180), CK => n50, RESET => n22, Q => Q(180)
                           );
   D_I_181 : FD_164 port map( D => d(181), CK => n50, RESET => n22, Q => Q(181)
                           );
   D_I_182 : FD_163 port map( D => d(182), CK => n50, RESET => n22, Q => Q(182)
                           );
   D_I_183 : FD_162 port map( D => d(183), CK => n50, RESET => n22, Q => Q(183)
                           );
   D_I_184 : FD_161 port map( D => d(184), CK => n50, RESET => n22, Q => Q(184)
                           );
   D_I_185 : FD_160 port map( D => d(185), CK => n50, RESET => n22, Q => Q(185)
                           );
   D_I_186 : FD_159 port map( D => d(186), CK => n50, RESET => n22, Q => Q(186)
                           );
   D_I_187 : FD_158 port map( D => d(187), CK => n51, RESET => n22, Q => Q(187)
                           );
   D_I_188 : FD_157 port map( D => d(188), CK => n51, RESET => n22, Q => Q(188)
                           );
   D_I_189 : FD_156 port map( D => d(189), CK => n51, RESET => n22, Q => Q(189)
                           );
   D_I_190 : FD_155 port map( D => d(190), CK => n51, RESET => n22, Q => Q(190)
                           );
   D_I_191 : FD_154 port map( D => d(191), CK => n51, RESET => n22, Q => Q(191)
                           );
   D_I_192 : FD_153 port map( D => d(192), CK => n51, RESET => n23, Q => Q(192)
                           );
   D_I_193 : FD_152 port map( D => d(193), CK => n51, RESET => n23, Q => Q(193)
                           );
   D_I_194 : FD_151 port map( D => d(194), CK => n51, RESET => n23, Q => Q(194)
                           );
   D_I_195 : FD_150 port map( D => d(195), CK => n51, RESET => n23, Q => Q(195)
                           );
   D_I_196 : FD_149 port map( D => d(196), CK => n51, RESET => n23, Q => Q(196)
                           );
   D_I_197 : FD_148 port map( D => d(197), CK => n51, RESET => n23, Q => Q(197)
                           );
   D_I_198 : FD_147 port map( D => d(198), CK => n52, RESET => n23, Q => Q(198)
                           );
   D_I_199 : FD_146 port map( D => d(199), CK => n52, RESET => n23, Q => Q(199)
                           );
   D_I_200 : FD_145 port map( D => d(200), CK => n52, RESET => n23, Q => Q(200)
                           );
   D_I_201 : FD_144 port map( D => d(201), CK => n52, RESET => n23, Q => Q(201)
                           );
   D_I_202 : FD_143 port map( D => d(202), CK => n52, RESET => n23, Q => Q(202)
                           );
   D_I_203 : FD_142 port map( D => d(203), CK => n52, RESET => n23, Q => Q(203)
                           );
   D_I_204 : FD_141 port map( D => d(204), CK => n52, RESET => n24, Q => Q(204)
                           );
   D_I_205 : FD_140 port map( D => d(205), CK => n52, RESET => n24, Q => Q(205)
                           );
   D_I_206 : FD_139 port map( D => d(206), CK => n52, RESET => n24, Q => Q(206)
                           );
   D_I_207 : FD_138 port map( D => d(207), CK => n52, RESET => n24, Q => Q(207)
                           );
   D_I_208 : FD_137 port map( D => d(208), CK => n52, RESET => n24, Q => Q(208)
                           );
   D_I_209 : FD_136 port map( D => d(209), CK => n53, RESET => n24, Q => Q(209)
                           );
   D_I_210 : FD_135 port map( D => d(210), CK => n53, RESET => n24, Q => Q(210)
                           );
   D_I_211 : FD_134 port map( D => d(211), CK => n53, RESET => n24, Q => Q(211)
                           );
   D_I_212 : FD_133 port map( D => d(212), CK => n53, RESET => n24, Q => Q(212)
                           );
   D_I_213 : FD_132 port map( D => d(213), CK => n53, RESET => n24, Q => Q(213)
                           );
   D_I_214 : FD_131 port map( D => d(214), CK => n53, RESET => n24, Q => Q(214)
                           );
   D_I_215 : FD_130 port map( D => d(215), CK => n53, RESET => n24, Q => Q(215)
                           );
   D_I_216 : FD_129 port map( D => d(216), CK => n53, RESET => n25, Q => Q(216)
                           );
   D_I_217 : FD_128 port map( D => d(217), CK => n53, RESET => n25, Q => Q(217)
                           );
   D_I_218 : FD_127 port map( D => d(218), CK => n53, RESET => n25, Q => Q(218)
                           );
   D_I_219 : FD_126 port map( D => d(219), CK => n53, RESET => n25, Q => Q(219)
                           );
   D_I_220 : FD_125 port map( D => d(220), CK => n54, RESET => n25, Q => Q(220)
                           );
   D_I_221 : FD_124 port map( D => d(221), CK => n54, RESET => n25, Q => Q(221)
                           );
   D_I_222 : FD_123 port map( D => d(222), CK => n54, RESET => n25, Q => Q(222)
                           );
   D_I_223 : FD_122 port map( D => d(223), CK => n54, RESET => n25, Q => Q(223)
                           );
   D_I_224 : FD_121 port map( D => d(224), CK => n54, RESET => n25, Q => Q(224)
                           );
   D_I_225 : FD_120 port map( D => d(225), CK => n54, RESET => n25, Q => Q(225)
                           );
   D_I_226 : FD_119 port map( D => d(226), CK => n54, RESET => n25, Q => Q(226)
                           );
   D_I_227 : FD_118 port map( D => d(227), CK => n54, RESET => n25, Q => Q(227)
                           );
   D_I_228 : FD_117 port map( D => d(228), CK => n54, RESET => n26, Q => Q(228)
                           );
   D_I_229 : FD_116 port map( D => d(229), CK => n54, RESET => n26, Q => Q(229)
                           );
   D_I_230 : FD_115 port map( D => d(230), CK => n54, RESET => n26, Q => Q(230)
                           );
   D_I_231 : FD_114 port map( D => d(231), CK => n55, RESET => n26, Q => Q(231)
                           );
   D_I_232 : FD_113 port map( D => d(232), CK => n55, RESET => n26, Q => Q(232)
                           );
   D_I_233 : FD_112 port map( D => d(233), CK => n55, RESET => n26, Q => Q(233)
                           );
   D_I_234 : FD_111 port map( D => d(234), CK => n55, RESET => n26, Q => Q(234)
                           );
   D_I_235 : FD_110 port map( D => d(235), CK => n55, RESET => n26, Q => Q(235)
                           );
   D_I_236 : FD_109 port map( D => d(236), CK => n55, RESET => n26, Q => Q(236)
                           );
   D_I_237 : FD_108 port map( D => d(237), CK => n55, RESET => n26, Q => Q(237)
                           );
   D_I_238 : FD_107 port map( D => d(238), CK => n55, RESET => n26, Q => Q(238)
                           );
   D_I_239 : FD_106 port map( D => d(239), CK => n55, RESET => n26, Q => Q(239)
                           );
   D_I_240 : FD_105 port map( D => d(240), CK => n55, RESET => n27, Q => Q(240)
                           );
   D_I_241 : FD_104 port map( D => d(241), CK => n55, RESET => n27, Q => Q(241)
                           );
   D_I_242 : FD_103 port map( D => d(242), CK => n56, RESET => n27, Q => Q(242)
                           );
   D_I_243 : FD_102 port map( D => d(243), CK => n56, RESET => n27, Q => Q(243)
                           );
   D_I_244 : FD_101 port map( D => d(244), CK => n56, RESET => n27, Q => Q(244)
                           );
   D_I_245 : FD_100 port map( D => d(245), CK => n56, RESET => n27, Q => Q(245)
                           );
   D_I_246 : FD_99 port map( D => d(246), CK => n56, RESET => n27, Q => Q(246))
                           ;
   D_I_247 : FD_98 port map( D => d(247), CK => n56, RESET => n27, Q => Q(247))
                           ;
   D_I_248 : FD_97 port map( D => d(248), CK => n56, RESET => n27, Q => Q(248))
                           ;
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_7 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_7;

architecture SYN_beh of encoder_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_6 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_6;

architecture SYN_beh of encoder_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_5 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_5;

architecture SYN_beh of encoder_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_4 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_4;

architecture SYN_beh of encoder_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_3 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_3;

architecture SYN_beh of encoder_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_2 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_2;

architecture SYN_beh of encoder_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_1 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_1;

architecture SYN_beh of encoder_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n33_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (32 downto 0);  Q 
         : out std_logic_vector (32 downto 0));

end reg_nbit_n33_1;

architecture SYN_struc of reg_nbit_n33_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1912
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1913
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1914
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1915
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1916
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1917
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1918
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1919
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1920
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1921
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1922
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1923
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1924
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1925
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1926
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1927
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1928
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1929
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1930
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1931
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1932
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1933
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1934
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1935
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1936
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1937
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1938
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1939
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1940
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1941
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1942
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1943
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1944
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1944 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1943 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1942 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1941 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1940 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1939 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1938 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1937 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1936 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1935 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1934 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1933 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1932 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1931 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1930 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1929 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1928 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1927 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1926 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1925 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1924 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1923 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1922 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1921 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1920 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1919 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1918 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1917 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1916 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1915 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1914 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1913 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   D_I_32 : FD_1912 port map( D => d(32), CK => n6, RESET => n3, Q => Q(32));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N32_Z1_4 is

   port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_zbit_nbit_N32_Z1_4;

architecture SYN_beh of MUX_zbit_nbit_N32_Z1_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n33, D => n7, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n33, D => n8, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n33, D => n9, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n33, D => n10, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n33, D => n11, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n33, D => n13, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n33, D => n14, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n33, D => n15, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n33, D => n16, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n33, D => n17, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n33, D => n18, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n33, D => n19, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n33, D => n20, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n33, D => n21, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n33, D => n22, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n33, D => n23, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n33, D => n24, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n33, D => n25, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n33, D => n26, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n33, D => n27, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n33, D => n28, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n33, D => n29, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n33, D => n30, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n33, D => n31, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n33, D => n32, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n33, D => n1, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n33, D => n2, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n33, D => n3, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n33, D => n4, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n33, D => n5, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n33, D => n6, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n33, D => n12, Q => Y(0));
   n33 <= '1';
   U3 : MUX2_X1 port map( A => inputs(25), B => inputs(57), S => SEL, Z => n1);
   U4 : MUX2_X1 port map( A => inputs(26), B => inputs(58), S => SEL, Z => n2);
   U5 : MUX2_X1 port map( A => inputs(27), B => inputs(59), S => SEL, Z => n3);
   U6 : MUX2_X1 port map( A => inputs(28), B => inputs(60), S => SEL, Z => n4);
   U7 : MUX2_X1 port map( A => inputs(29), B => inputs(61), S => SEL, Z => n5);
   U8 : MUX2_X1 port map( A => inputs(30), B => inputs(62), S => SEL, Z => n6);
   U9 : MUX2_X1 port map( A => inputs(0), B => inputs(32), S => SEL, Z => n7);
   U10 : MUX2_X1 port map( A => inputs(1), B => inputs(33), S => SEL, Z => n8);
   U11 : MUX2_X1 port map( A => inputs(2), B => inputs(34), S => SEL, Z => n9);
   U12 : MUX2_X1 port map( A => inputs(3), B => inputs(35), S => SEL, Z => n10)
                           ;
   U13 : MUX2_X1 port map( A => inputs(4), B => inputs(36), S => SEL, Z => n11)
                           ;
   U14 : MUX2_X1 port map( A => inputs(31), B => inputs(63), S => SEL, Z => n12
                           );
   U15 : MUX2_X1 port map( A => inputs(5), B => inputs(37), S => SEL, Z => n13)
                           ;
   U16 : MUX2_X1 port map( A => inputs(6), B => inputs(38), S => SEL, Z => n14)
                           ;
   U17 : MUX2_X1 port map( A => inputs(7), B => inputs(39), S => SEL, Z => n15)
                           ;
   U18 : MUX2_X1 port map( A => inputs(8), B => inputs(40), S => SEL, Z => n16)
                           ;
   U19 : MUX2_X1 port map( A => inputs(9), B => inputs(41), S => SEL, Z => n17)
                           ;
   U20 : MUX2_X1 port map( A => inputs(10), B => inputs(42), S => SEL, Z => n18
                           );
   U21 : MUX2_X1 port map( A => inputs(11), B => inputs(43), S => SEL, Z => n19
                           );
   U22 : MUX2_X1 port map( A => inputs(12), B => inputs(44), S => SEL, Z => n20
                           );
   U23 : MUX2_X1 port map( A => inputs(13), B => inputs(45), S => SEL, Z => n21
                           );
   U24 : MUX2_X1 port map( A => inputs(14), B => inputs(46), S => SEL, Z => n22
                           );
   U25 : MUX2_X1 port map( A => inputs(15), B => inputs(47), S => SEL, Z => n23
                           );
   U26 : MUX2_X1 port map( A => inputs(16), B => inputs(48), S => SEL, Z => n24
                           );
   U27 : MUX2_X1 port map( A => inputs(17), B => inputs(49), S => SEL, Z => n25
                           );
   U28 : MUX2_X1 port map( A => inputs(18), B => inputs(50), S => SEL, Z => n26
                           );
   U29 : MUX2_X1 port map( A => inputs(19), B => inputs(51), S => SEL, Z => n27
                           );
   U30 : MUX2_X1 port map( A => inputs(20), B => inputs(52), S => SEL, Z => n28
                           );
   U31 : MUX2_X1 port map( A => inputs(21), B => inputs(53), S => SEL, Z => n29
                           );
   U32 : MUX2_X1 port map( A => inputs(22), B => inputs(54), S => SEL, Z => n30
                           );
   U33 : MUX2_X1 port map( A => inputs(23), B => inputs(55), S => SEL, Z => n31
                           );
   U34 : MUX2_X1 port map( A => inputs(24), B => inputs(56), S => SEL, Z => n32
                           );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N32_Z1_3 is

   port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_zbit_nbit_N32_Z1_3;

architecture SYN_beh of MUX_zbit_nbit_N32_Z1_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n33, D => n7, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n33, D => n8, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n33, D => n9, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n33, D => n10, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n33, D => n11, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n33, D => n13, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n33, D => n14, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n33, D => n15, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n33, D => n16, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n33, D => n17, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n33, D => n18, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n33, D => n19, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n33, D => n20, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n33, D => n21, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n33, D => n22, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n33, D => n23, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n33, D => n24, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n33, D => n25, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n33, D => n26, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n33, D => n27, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n33, D => n28, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n33, D => n29, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n33, D => n30, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n33, D => n31, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n33, D => n32, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n33, D => n1, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n33, D => n2, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n33, D => n3, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n33, D => n4, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n33, D => n5, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n33, D => n6, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n33, D => n12, Q => Y(0));
   n33 <= '1';
   U3 : MUX2_X1 port map( A => inputs(25), B => inputs(57), S => SEL, Z => n1);
   U4 : MUX2_X1 port map( A => inputs(26), B => inputs(58), S => SEL, Z => n2);
   U5 : MUX2_X1 port map( A => inputs(27), B => inputs(59), S => SEL, Z => n3);
   U6 : MUX2_X1 port map( A => inputs(28), B => inputs(60), S => SEL, Z => n4);
   U7 : MUX2_X1 port map( A => inputs(29), B => inputs(61), S => SEL, Z => n5);
   U8 : MUX2_X1 port map( A => inputs(30), B => inputs(62), S => SEL, Z => n6);
   U9 : MUX2_X1 port map( A => inputs(0), B => inputs(32), S => SEL, Z => n7);
   U10 : MUX2_X1 port map( A => inputs(1), B => inputs(33), S => SEL, Z => n8);
   U11 : MUX2_X1 port map( A => inputs(2), B => inputs(34), S => SEL, Z => n9);
   U12 : MUX2_X1 port map( A => inputs(3), B => inputs(35), S => SEL, Z => n10)
                           ;
   U13 : MUX2_X1 port map( A => inputs(4), B => inputs(36), S => SEL, Z => n11)
                           ;
   U14 : MUX2_X1 port map( A => inputs(31), B => inputs(63), S => SEL, Z => n12
                           );
   U15 : MUX2_X1 port map( A => inputs(5), B => inputs(37), S => SEL, Z => n13)
                           ;
   U16 : MUX2_X1 port map( A => inputs(6), B => inputs(38), S => SEL, Z => n14)
                           ;
   U17 : MUX2_X1 port map( A => inputs(7), B => inputs(39), S => SEL, Z => n15)
                           ;
   U18 : MUX2_X1 port map( A => inputs(8), B => inputs(40), S => SEL, Z => n16)
                           ;
   U19 : MUX2_X1 port map( A => inputs(9), B => inputs(41), S => SEL, Z => n17)
                           ;
   U20 : MUX2_X1 port map( A => inputs(10), B => inputs(42), S => SEL, Z => n18
                           );
   U21 : MUX2_X1 port map( A => inputs(11), B => inputs(43), S => SEL, Z => n19
                           );
   U22 : MUX2_X1 port map( A => inputs(12), B => inputs(44), S => SEL, Z => n20
                           );
   U23 : MUX2_X1 port map( A => inputs(13), B => inputs(45), S => SEL, Z => n21
                           );
   U24 : MUX2_X1 port map( A => inputs(14), B => inputs(46), S => SEL, Z => n22
                           );
   U25 : MUX2_X1 port map( A => inputs(15), B => inputs(47), S => SEL, Z => n23
                           );
   U26 : MUX2_X1 port map( A => inputs(16), B => inputs(48), S => SEL, Z => n24
                           );
   U27 : MUX2_X1 port map( A => inputs(17), B => inputs(49), S => SEL, Z => n25
                           );
   U28 : MUX2_X1 port map( A => inputs(18), B => inputs(50), S => SEL, Z => n26
                           );
   U29 : MUX2_X1 port map( A => inputs(19), B => inputs(51), S => SEL, Z => n27
                           );
   U30 : MUX2_X1 port map( A => inputs(20), B => inputs(52), S => SEL, Z => n28
                           );
   U31 : MUX2_X1 port map( A => inputs(21), B => inputs(53), S => SEL, Z => n29
                           );
   U32 : MUX2_X1 port map( A => inputs(22), B => inputs(54), S => SEL, Z => n30
                           );
   U33 : MUX2_X1 port map( A => inputs(23), B => inputs(55), S => SEL, Z => n31
                           );
   U34 : MUX2_X1 port map( A => inputs(24), B => inputs(56), S => SEL, Z => n32
                           );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N32_Z1_2 is

   port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_zbit_nbit_N32_Z1_2;

architecture SYN_beh of MUX_zbit_nbit_N32_Z1_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n33, D => n32, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n33, D => n31, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n33, D => n30, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n33, D => n29, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n33, D => n28, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n33, D => n27, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n33, D => n26, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n33, D => n25, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n33, D => n24, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n33, D => n23, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n33, D => n22, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n33, D => n21, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n33, D => n20, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n33, D => n19, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n33, D => n18, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n33, D => n17, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n33, D => n16, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n33, D => n15, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n33, D => n14, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n33, D => n13, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n33, D => n12, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n33, D => n11, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n33, D => n10, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n33, D => n9, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n33, D => n8, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n33, D => n7, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n33, D => n6, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n33, D => n5, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n33, D => n4, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n33, D => n3, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n33, D => n2, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n33, D => n1, Q => Y(0));
   n33 <= '1';
   U3 : MUX2_X1 port map( A => inputs(31), B => inputs(63), S => SEL, Z => n1);
   U4 : MUX2_X1 port map( A => inputs(30), B => inputs(62), S => SEL, Z => n2);
   U5 : MUX2_X1 port map( A => inputs(29), B => inputs(61), S => SEL, Z => n3);
   U6 : MUX2_X1 port map( A => inputs(28), B => inputs(60), S => SEL, Z => n4);
   U7 : MUX2_X1 port map( A => inputs(27), B => inputs(59), S => SEL, Z => n5);
   U8 : MUX2_X1 port map( A => inputs(26), B => inputs(58), S => SEL, Z => n6);
   U9 : MUX2_X1 port map( A => inputs(25), B => inputs(57), S => SEL, Z => n7);
   U10 : MUX2_X1 port map( A => inputs(24), B => inputs(56), S => SEL, Z => n8)
                           ;
   U11 : MUX2_X1 port map( A => inputs(23), B => inputs(55), S => SEL, Z => n9)
                           ;
   U12 : MUX2_X1 port map( A => inputs(22), B => inputs(54), S => SEL, Z => n10
                           );
   U13 : MUX2_X1 port map( A => inputs(21), B => inputs(53), S => SEL, Z => n11
                           );
   U14 : MUX2_X1 port map( A => inputs(20), B => inputs(52), S => SEL, Z => n12
                           );
   U15 : MUX2_X1 port map( A => inputs(19), B => inputs(51), S => SEL, Z => n13
                           );
   U16 : MUX2_X1 port map( A => inputs(18), B => inputs(50), S => SEL, Z => n14
                           );
   U17 : MUX2_X1 port map( A => inputs(17), B => inputs(49), S => SEL, Z => n15
                           );
   U18 : MUX2_X1 port map( A => inputs(16), B => inputs(48), S => SEL, Z => n16
                           );
   U19 : MUX2_X1 port map( A => inputs(15), B => inputs(47), S => SEL, Z => n17
                           );
   U20 : MUX2_X1 port map( A => inputs(14), B => inputs(46), S => SEL, Z => n18
                           );
   U21 : MUX2_X1 port map( A => inputs(13), B => inputs(45), S => SEL, Z => n19
                           );
   U22 : MUX2_X1 port map( A => inputs(12), B => inputs(44), S => SEL, Z => n20
                           );
   U23 : MUX2_X1 port map( A => inputs(11), B => inputs(43), S => SEL, Z => n21
                           );
   U24 : MUX2_X1 port map( A => inputs(10), B => inputs(42), S => SEL, Z => n22
                           );
   U25 : MUX2_X1 port map( A => inputs(9), B => inputs(41), S => SEL, Z => n23)
                           ;
   U26 : MUX2_X1 port map( A => inputs(8), B => inputs(40), S => SEL, Z => n24)
                           ;
   U27 : MUX2_X1 port map( A => inputs(7), B => inputs(39), S => SEL, Z => n25)
                           ;
   U28 : MUX2_X1 port map( A => inputs(6), B => inputs(38), S => SEL, Z => n26)
                           ;
   U29 : MUX2_X1 port map( A => inputs(5), B => inputs(37), S => SEL, Z => n27)
                           ;
   U30 : MUX2_X1 port map( A => inputs(4), B => inputs(36), S => SEL, Z => n28)
                           ;
   U31 : MUX2_X1 port map( A => inputs(3), B => inputs(35), S => SEL, Z => n29)
                           ;
   U32 : MUX2_X1 port map( A => inputs(2), B => inputs(34), S => SEL, Z => n30)
                           ;
   U33 : MUX2_X1 port map( A => inputs(1), B => inputs(33), S => SEL, Z => n31)
                           ;
   U34 : MUX2_X1 port map( A => inputs(0), B => inputs(32), S => SEL, Z => n32)
                           ;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N32_Z1_1 is

   port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_zbit_nbit_N32_Z1_1;

architecture SYN_beh of MUX_zbit_nbit_N32_Z1_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n33, D => n7, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n33, D => n8, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n33, D => n9, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n33, D => n10, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n33, D => n11, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n33, D => n13, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n33, D => n14, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n33, D => n15, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n33, D => n16, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n33, D => n17, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n33, D => n18, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n33, D => n19, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n33, D => n20, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n33, D => n21, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n33, D => n22, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n33, D => n23, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n33, D => n24, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n33, D => n25, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n33, D => n26, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n33, D => n27, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n33, D => n28, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n33, D => n29, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n33, D => n30, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n33, D => n31, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n33, D => n32, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n33, D => n1, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n33, D => n2, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n33, D => n3, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n33, D => n4, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n33, D => n5, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n33, D => n6, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n33, D => n12, Q => Y(0));
   n33 <= '1';
   U3 : MUX2_X1 port map( A => inputs(25), B => inputs(57), S => SEL, Z => n1);
   U4 : MUX2_X1 port map( A => inputs(26), B => inputs(58), S => SEL, Z => n2);
   U5 : MUX2_X1 port map( A => inputs(27), B => inputs(59), S => SEL, Z => n3);
   U6 : MUX2_X1 port map( A => inputs(28), B => inputs(60), S => SEL, Z => n4);
   U7 : MUX2_X1 port map( A => inputs(29), B => inputs(61), S => SEL, Z => n5);
   U8 : MUX2_X1 port map( A => inputs(30), B => inputs(62), S => SEL, Z => n6);
   U9 : MUX2_X1 port map( A => inputs(0), B => inputs(32), S => SEL, Z => n7);
   U10 : MUX2_X1 port map( A => inputs(1), B => inputs(33), S => SEL, Z => n8);
   U11 : MUX2_X1 port map( A => inputs(2), B => inputs(34), S => SEL, Z => n9);
   U12 : MUX2_X1 port map( A => inputs(3), B => inputs(35), S => SEL, Z => n10)
                           ;
   U13 : MUX2_X1 port map( A => inputs(4), B => inputs(36), S => SEL, Z => n11)
                           ;
   U14 : MUX2_X1 port map( A => inputs(31), B => inputs(63), S => SEL, Z => n12
                           );
   U15 : MUX2_X1 port map( A => inputs(5), B => inputs(37), S => SEL, Z => n13)
                           ;
   U16 : MUX2_X1 port map( A => inputs(6), B => inputs(38), S => SEL, Z => n14)
                           ;
   U17 : MUX2_X1 port map( A => inputs(7), B => inputs(39), S => SEL, Z => n15)
                           ;
   U18 : MUX2_X1 port map( A => inputs(8), B => inputs(40), S => SEL, Z => n16)
                           ;
   U19 : MUX2_X1 port map( A => inputs(9), B => inputs(41), S => SEL, Z => n17)
                           ;
   U20 : MUX2_X1 port map( A => inputs(10), B => inputs(42), S => SEL, Z => n18
                           );
   U21 : MUX2_X1 port map( A => inputs(11), B => inputs(43), S => SEL, Z => n19
                           );
   U22 : MUX2_X1 port map( A => inputs(12), B => inputs(44), S => SEL, Z => n20
                           );
   U23 : MUX2_X1 port map( A => inputs(13), B => inputs(45), S => SEL, Z => n21
                           );
   U24 : MUX2_X1 port map( A => inputs(14), B => inputs(46), S => SEL, Z => n22
                           );
   U25 : MUX2_X1 port map( A => inputs(15), B => inputs(47), S => SEL, Z => n23
                           );
   U26 : MUX2_X1 port map( A => inputs(16), B => inputs(48), S => SEL, Z => n24
                           );
   U27 : MUX2_X1 port map( A => inputs(17), B => inputs(49), S => SEL, Z => n25
                           );
   U28 : MUX2_X1 port map( A => inputs(18), B => inputs(50), S => SEL, Z => n26
                           );
   U29 : MUX2_X1 port map( A => inputs(19), B => inputs(51), S => SEL, Z => n27
                           );
   U30 : MUX2_X1 port map( A => inputs(20), B => inputs(52), S => SEL, Z => n28
                           );
   U31 : MUX2_X1 port map( A => inputs(21), B => inputs(53), S => SEL, Z => n29
                           );
   U32 : MUX2_X1 port map( A => inputs(22), B => inputs(54), S => SEL, Z => n30
                           );
   U33 : MUX2_X1 port map( A => inputs(23), B => inputs(55), S => SEL, Z => n31
                           );
   U34 : MUX2_X1 port map( A => inputs(24), B => inputs(56), S => SEL, Z => n32
                           );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n5_2 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  Q :
         out std_logic_vector (4 downto 0));

end reg_nbit_n5_2;

architecture SYN_struc of reg_nbit_n5_2 is

   component FD_2079
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2080
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2081
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2082
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2083
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;

begin
   
   D_I_0 : FD_2083 port map( D => d(0), CK => clk, RESET => reset, Q => Q(0));
   D_I_1 : FD_2082 port map( D => d(1), CK => clk, RESET => reset, Q => Q(1));
   D_I_2 : FD_2081 port map( D => d(2), CK => clk, RESET => reset, Q => Q(2));
   D_I_3 : FD_2080 port map( D => d(3), CK => clk, RESET => reset, Q => Q(3));
   D_I_4 : FD_2079 port map( D => d(4), CK => clk, RESET => reset, Q => Q(4));

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n5_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  Q :
         out std_logic_vector (4 downto 0));

end reg_nbit_n5_1;

architecture SYN_struc of reg_nbit_n5_1 is

   component FD_2074
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2075
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2076
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2077
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2078
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;

begin
   
   D_I_0 : FD_2078 port map( D => d(0), CK => clk, RESET => reset, Q => Q(0));
   D_I_1 : FD_2077 port map( D => d(1), CK => clk, RESET => reset, Q => Q(1));
   D_I_2 : FD_2076 port map( D => d(2), CK => clk, RESET => reset, Q => Q(2));
   D_I_3 : FD_2075 port map( D => d(3), CK => clk, RESET => reset, Q => Q(3));
   D_I_4 : FD_2074 port map( D => d(4), CK => clk, RESET => reset, Q => Q(4));

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_15 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_15;

architecture SYN_struc of reg_nbit_n32_15 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2121
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2122
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2123
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2124
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2125
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2126
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2127
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2128
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2129
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2130
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2131
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2132
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2133
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2134
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2135
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2136
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2137
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2138
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2139
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2140
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2141
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2142
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2143
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2144
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2145
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2146
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2147
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2148
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2149
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2150
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2151
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2152
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_2152 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_2151 port map( D => d(1), CK => n1, RESET => reset, Q => Q(1));
   D_I_2 : FD_2150 port map( D => d(2), CK => n1, RESET => reset, Q => Q(2));
   D_I_3 : FD_2149 port map( D => d(3), CK => n1, RESET => reset, Q => Q(3));
   D_I_4 : FD_2148 port map( D => d(4), CK => n1, RESET => reset, Q => Q(4));
   D_I_5 : FD_2147 port map( D => d(5), CK => n1, RESET => reset, Q => Q(5));
   D_I_6 : FD_2146 port map( D => d(6), CK => n1, RESET => reset, Q => Q(6));
   D_I_7 : FD_2145 port map( D => d(7), CK => n1, RESET => reset, Q => Q(7));
   D_I_8 : FD_2144 port map( D => d(8), CK => n1, RESET => reset, Q => Q(8));
   D_I_9 : FD_2143 port map( D => d(9), CK => n1, RESET => reset, Q => Q(9));
   D_I_10 : FD_2142 port map( D => d(10), CK => n1, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2141 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2140 port map( D => d(12), CK => n2, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2139 port map( D => d(13), CK => n2, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2138 port map( D => d(14), CK => n2, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2137 port map( D => d(15), CK => n2, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2136 port map( D => d(16), CK => n2, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2135 port map( D => d(17), CK => n2, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2134 port map( D => d(18), CK => n2, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2133 port map( D => d(19), CK => n2, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2132 port map( D => d(20), CK => n2, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2131 port map( D => d(21), CK => n2, RESET => reset, Q => Q(21))
                           ;
   D_I_22 : FD_2130 port map( D => d(22), CK => n3, RESET => reset, Q => Q(22))
                           ;
   D_I_23 : FD_2129 port map( D => d(23), CK => n3, RESET => reset, Q => Q(23))
                           ;
   D_I_24 : FD_2128 port map( D => d(24), CK => n3, RESET => reset, Q => Q(24))
                           ;
   D_I_25 : FD_2127 port map( D => d(25), CK => n3, RESET => reset, Q => Q(25))
                           ;
   D_I_26 : FD_2126 port map( D => d(26), CK => n3, RESET => reset, Q => Q(26))
                           ;
   D_I_27 : FD_2125 port map( D => d(27), CK => n3, RESET => reset, Q => Q(27))
                           ;
   D_I_28 : FD_2124 port map( D => d(28), CK => n3, RESET => reset, Q => Q(28))
                           ;
   D_I_29 : FD_2123 port map( D => d(29), CK => n3, RESET => reset, Q => Q(29))
                           ;
   D_I_30 : FD_2122 port map( D => d(30), CK => n3, RESET => reset, Q => Q(30))
                           ;
   D_I_31 : FD_2121 port map( D => d(31), CK => n3, RESET => reset, Q => Q(31))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n1);
   U2 : BUF_X1 port map( A => clk, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_14 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_14;

architecture SYN_struc of reg_nbit_n32_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2089
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2090
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2091
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2092
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2093
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2094
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2095
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2096
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2097
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2098
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2099
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2100
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2101
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2102
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2103
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2104
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2105
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2106
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2107
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2108
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2109
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2110
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2111
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2112
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2113
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2114
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2115
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2116
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2117
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2118
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2119
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2120
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_2120 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_2119 port map( D => d(1), CK => n1, RESET => reset, Q => Q(1));
   D_I_2 : FD_2118 port map( D => d(2), CK => n1, RESET => reset, Q => Q(2));
   D_I_3 : FD_2117 port map( D => d(3), CK => n1, RESET => reset, Q => Q(3));
   D_I_4 : FD_2116 port map( D => d(4), CK => n1, RESET => reset, Q => Q(4));
   D_I_5 : FD_2115 port map( D => d(5), CK => n1, RESET => reset, Q => Q(5));
   D_I_6 : FD_2114 port map( D => d(6), CK => n1, RESET => reset, Q => Q(6));
   D_I_7 : FD_2113 port map( D => d(7), CK => n1, RESET => reset, Q => Q(7));
   D_I_8 : FD_2112 port map( D => d(8), CK => n1, RESET => reset, Q => Q(8));
   D_I_9 : FD_2111 port map( D => d(9), CK => n1, RESET => reset, Q => Q(9));
   D_I_10 : FD_2110 port map( D => d(10), CK => n1, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2109 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2108 port map( D => d(12), CK => n2, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2107 port map( D => d(13), CK => n2, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2106 port map( D => d(14), CK => n2, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2105 port map( D => d(15), CK => n2, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2104 port map( D => d(16), CK => n2, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2103 port map( D => d(17), CK => n2, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2102 port map( D => d(18), CK => n2, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2101 port map( D => d(19), CK => n2, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2100 port map( D => d(20), CK => n2, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2099 port map( D => d(21), CK => n2, RESET => reset, Q => Q(21))
                           ;
   D_I_22 : FD_2098 port map( D => d(22), CK => n3, RESET => reset, Q => Q(22))
                           ;
   D_I_23 : FD_2097 port map( D => d(23), CK => n3, RESET => reset, Q => Q(23))
                           ;
   D_I_24 : FD_2096 port map( D => d(24), CK => n3, RESET => reset, Q => Q(24))
                           ;
   D_I_25 : FD_2095 port map( D => d(25), CK => n3, RESET => reset, Q => Q(25))
                           ;
   D_I_26 : FD_2094 port map( D => d(26), CK => n3, RESET => reset, Q => Q(26))
                           ;
   D_I_27 : FD_2093 port map( D => d(27), CK => n3, RESET => reset, Q => Q(27))
                           ;
   D_I_28 : FD_2092 port map( D => d(28), CK => n3, RESET => reset, Q => Q(28))
                           ;
   D_I_29 : FD_2091 port map( D => d(29), CK => n3, RESET => reset, Q => Q(29))
                           ;
   D_I_30 : FD_2090 port map( D => d(30), CK => n3, RESET => reset, Q => Q(30))
                           ;
   D_I_31 : FD_2089 port map( D => d(31), CK => n3, RESET => reset, Q => Q(31))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n1);
   U2 : BUF_X1 port map( A => clk, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_13 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_13;

architecture SYN_struc of reg_nbit_n32_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2042
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2043
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2044
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2045
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2046
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2047
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2048
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2049
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2050
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2051
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2052
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2053
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2054
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2055
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2056
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2057
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2058
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2059
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2060
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2061
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2062
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2063
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2064
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2065
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2066
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2067
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2068
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2069
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2070
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2071
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2072
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2073
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_2073 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_2072 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_2071 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_2070 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_2069 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_2068 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_2067 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_2066 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_2065 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_2064 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_2063 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_2062 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_2061 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_2060 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_2059 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_2058 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_2057 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_2056 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_2055 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_2054 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_2053 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_2052 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_2051 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_2050 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_2049 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_2048 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_2047 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_2046 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_2045 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_2044 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_2043 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_2042 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_12 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_12;

architecture SYN_struc of reg_nbit_n32_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2010
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2011
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2012
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2013
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2014
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2015
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2016
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2017
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2018
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2019
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2020
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2021
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2022
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2023
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2024
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2025
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2026
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2027
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2028
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2029
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2030
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2031
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2032
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2033
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2034
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2035
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2036
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2037
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2038
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2039
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2040
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2041
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_2041 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_2040 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_2039 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_2038 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_2037 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_2036 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_2035 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_2034 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_2033 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_2032 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_2031 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_2030 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_2029 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_2028 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_2027 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_2026 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_2025 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_2024 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_2023 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_2022 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_2021 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_2020 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_2019 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_2018 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_2017 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_2016 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_2015 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_2014 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_2013 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_2012 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_2011 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_2010 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_11 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_11;

architecture SYN_struc of reg_nbit_n32_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1978
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1979
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1980
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1981
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1982
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1983
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1984
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1985
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1986
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1987
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1988
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1989
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1990
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1991
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1992
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1993
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1994
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1995
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1996
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1997
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1998
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1999
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2000
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2001
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2002
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2003
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2004
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2005
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2006
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2007
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2008
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2009
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_2009 port map( D => d(0), CK => clk, RESET => n1, Q => Q(0));
   D_I_1 : FD_2008 port map( D => d(1), CK => clk, RESET => n1, Q => Q(1));
   D_I_2 : FD_2007 port map( D => d(2), CK => clk, RESET => n1, Q => Q(2));
   D_I_3 : FD_2006 port map( D => d(3), CK => clk, RESET => n1, Q => Q(3));
   D_I_4 : FD_2005 port map( D => d(4), CK => clk, RESET => n1, Q => Q(4));
   D_I_5 : FD_2004 port map( D => d(5), CK => clk, RESET => n1, Q => Q(5));
   D_I_6 : FD_2003 port map( D => d(6), CK => clk, RESET => n1, Q => Q(6));
   D_I_7 : FD_2002 port map( D => d(7), CK => clk, RESET => n1, Q => Q(7));
   D_I_8 : FD_2001 port map( D => d(8), CK => clk, RESET => n1, Q => Q(8));
   D_I_9 : FD_2000 port map( D => d(9), CK => clk, RESET => n1, Q => Q(9));
   D_I_10 : FD_1999 port map( D => d(10), CK => clk, RESET => n1, Q => Q(10));
   D_I_11 : FD_1998 port map( D => d(11), CK => clk, RESET => n1, Q => Q(11));
   D_I_12 : FD_1997 port map( D => d(12), CK => clk, RESET => n2, Q => Q(12));
   D_I_13 : FD_1996 port map( D => d(13), CK => clk, RESET => n2, Q => Q(13));
   D_I_14 : FD_1995 port map( D => d(14), CK => clk, RESET => n2, Q => Q(14));
   D_I_15 : FD_1994 port map( D => d(15), CK => clk, RESET => n2, Q => Q(15));
   D_I_16 : FD_1993 port map( D => d(16), CK => clk, RESET => n2, Q => Q(16));
   D_I_17 : FD_1992 port map( D => d(17), CK => clk, RESET => n2, Q => Q(17));
   D_I_18 : FD_1991 port map( D => d(18), CK => clk, RESET => n2, Q => Q(18));
   D_I_19 : FD_1990 port map( D => d(19), CK => clk, RESET => n2, Q => Q(19));
   D_I_20 : FD_1989 port map( D => d(20), CK => clk, RESET => n2, Q => Q(20));
   D_I_21 : FD_1988 port map( D => d(21), CK => clk, RESET => n2, Q => Q(21));
   D_I_22 : FD_1987 port map( D => d(22), CK => clk, RESET => n2, Q => Q(22));
   D_I_23 : FD_1986 port map( D => d(23), CK => clk, RESET => n2, Q => Q(23));
   D_I_24 : FD_1985 port map( D => d(24), CK => clk, RESET => n3, Q => Q(24));
   D_I_25 : FD_1984 port map( D => d(25), CK => clk, RESET => n3, Q => Q(25));
   D_I_26 : FD_1983 port map( D => d(26), CK => clk, RESET => n3, Q => Q(26));
   D_I_27 : FD_1982 port map( D => d(27), CK => clk, RESET => n3, Q => Q(27));
   D_I_28 : FD_1981 port map( D => d(28), CK => clk, RESET => n3, Q => Q(28));
   D_I_29 : FD_1980 port map( D => d(29), CK => clk, RESET => n3, Q => Q(29));
   D_I_30 : FD_1979 port map( D => d(30), CK => clk, RESET => n3, Q => Q(30));
   D_I_31 : FD_1978 port map( D => d(31), CK => clk, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_10 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_10;

architecture SYN_struc of reg_nbit_n32_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1879
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1880
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1881
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1882
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1883
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1884
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1885
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1886
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1887
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1888
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1889
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1890
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1891
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1892
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1893
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1894
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1895
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1896
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1897
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1898
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1899
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1900
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1901
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1902
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1903
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1904
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1905
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1906
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1907
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1908
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1909
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1910
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1910 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1909 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1908 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1907 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1906 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1905 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1904 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1903 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1902 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1901 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1900 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1899 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1898 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1897 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1896 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1895 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1894 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1893 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1892 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1891 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1890 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1889 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1888 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1887 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1886 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1885 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1884 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1883 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1882 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1881 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1880 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1879 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_9 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_9;

architecture SYN_struc of reg_nbit_n32_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1847
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1848
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1849
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1850
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1851
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1852
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1853
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1854
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1855
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1856
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1857
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1858
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1859
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1860
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1861
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1862
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1863
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1864
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1865
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1866
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1867
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1868
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1869
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1870
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1871
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1872
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1873
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1874
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1875
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1876
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1877
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1878
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1878 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1877 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1876 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1875 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1874 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1873 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1872 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1871 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1870 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1869 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1868 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1867 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1866 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1865 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1864 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1863 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1862 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1861 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1860 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1859 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1858 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1857 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1856 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1855 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1854 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1853 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1852 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1851 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1850 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1849 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1848 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1847 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_8 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_8;

architecture SYN_struc of reg_nbit_n32_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1815
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1816
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1817
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1818
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1819
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1820
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1821
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1822
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1823
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1824
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1825
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1826
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1827
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1828
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1829
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1830
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1831
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1832
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1833
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1834
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1835
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1836
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1837
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1838
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1839
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1840
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1841
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1842
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1843
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1844
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1845
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1846
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_1846 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_1845 port map( D => d(1), CK => n1, RESET => reset, Q => Q(1));
   D_I_2 : FD_1844 port map( D => d(2), CK => n1, RESET => reset, Q => Q(2));
   D_I_3 : FD_1843 port map( D => d(3), CK => n1, RESET => reset, Q => Q(3));
   D_I_4 : FD_1842 port map( D => d(4), CK => n1, RESET => reset, Q => Q(4));
   D_I_5 : FD_1841 port map( D => d(5), CK => n1, RESET => reset, Q => Q(5));
   D_I_6 : FD_1840 port map( D => d(6), CK => n1, RESET => reset, Q => Q(6));
   D_I_7 : FD_1839 port map( D => d(7), CK => n1, RESET => reset, Q => Q(7));
   D_I_8 : FD_1838 port map( D => d(8), CK => n1, RESET => reset, Q => Q(8));
   D_I_9 : FD_1837 port map( D => d(9), CK => n1, RESET => reset, Q => Q(9));
   D_I_10 : FD_1836 port map( D => d(10), CK => n1, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_1835 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_1834 port map( D => d(12), CK => n2, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_1833 port map( D => d(13), CK => n2, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_1832 port map( D => d(14), CK => n2, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_1831 port map( D => d(15), CK => n2, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_1830 port map( D => d(16), CK => n2, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_1829 port map( D => d(17), CK => n2, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_1828 port map( D => d(18), CK => n2, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_1827 port map( D => d(19), CK => n2, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_1826 port map( D => d(20), CK => n2, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_1825 port map( D => d(21), CK => n2, RESET => reset, Q => Q(21))
                           ;
   D_I_22 : FD_1824 port map( D => d(22), CK => n3, RESET => reset, Q => Q(22))
                           ;
   D_I_23 : FD_1823 port map( D => d(23), CK => n3, RESET => reset, Q => Q(23))
                           ;
   D_I_24 : FD_1822 port map( D => d(24), CK => n3, RESET => reset, Q => Q(24))
                           ;
   D_I_25 : FD_1821 port map( D => d(25), CK => n3, RESET => reset, Q => Q(25))
                           ;
   D_I_26 : FD_1820 port map( D => d(26), CK => n3, RESET => reset, Q => Q(26))
                           ;
   D_I_27 : FD_1819 port map( D => d(27), CK => n3, RESET => reset, Q => Q(27))
                           ;
   D_I_28 : FD_1818 port map( D => d(28), CK => n3, RESET => reset, Q => Q(28))
                           ;
   D_I_29 : FD_1817 port map( D => d(29), CK => n3, RESET => reset, Q => Q(29))
                           ;
   D_I_30 : FD_1816 port map( D => d(30), CK => n3, RESET => reset, Q => Q(30))
                           ;
   D_I_31 : FD_1815 port map( D => d(31), CK => n3, RESET => reset, Q => Q(31))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n1);
   U2 : BUF_X1 port map( A => clk, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_7 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_7;

architecture SYN_struc of reg_nbit_n32_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1783
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1784
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1785
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1786
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1787
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1788
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1789
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1790
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1791
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1792
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1793
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1794
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1795
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1796
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1797
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1798
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1799
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1800
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1801
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1802
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1803
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1804
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1805
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1806
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1807
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1808
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1809
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1810
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1811
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1812
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1813
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1814
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_1814 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_1813 port map( D => d(1), CK => n1, RESET => reset, Q => Q(1));
   D_I_2 : FD_1812 port map( D => d(2), CK => n1, RESET => reset, Q => Q(2));
   D_I_3 : FD_1811 port map( D => d(3), CK => n1, RESET => reset, Q => Q(3));
   D_I_4 : FD_1810 port map( D => d(4), CK => n1, RESET => reset, Q => Q(4));
   D_I_5 : FD_1809 port map( D => d(5), CK => n1, RESET => reset, Q => Q(5));
   D_I_6 : FD_1808 port map( D => d(6), CK => n1, RESET => reset, Q => Q(6));
   D_I_7 : FD_1807 port map( D => d(7), CK => n1, RESET => reset, Q => Q(7));
   D_I_8 : FD_1806 port map( D => d(8), CK => n1, RESET => reset, Q => Q(8));
   D_I_9 : FD_1805 port map( D => d(9), CK => n1, RESET => reset, Q => Q(9));
   D_I_10 : FD_1804 port map( D => d(10), CK => n1, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_1803 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_1802 port map( D => d(12), CK => n2, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_1801 port map( D => d(13), CK => n2, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_1800 port map( D => d(14), CK => n2, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_1799 port map( D => d(15), CK => n2, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_1798 port map( D => d(16), CK => n2, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_1797 port map( D => d(17), CK => n2, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_1796 port map( D => d(18), CK => n2, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_1795 port map( D => d(19), CK => n2, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_1794 port map( D => d(20), CK => n2, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_1793 port map( D => d(21), CK => n2, RESET => reset, Q => Q(21))
                           ;
   D_I_22 : FD_1792 port map( D => d(22), CK => n3, RESET => reset, Q => Q(22))
                           ;
   D_I_23 : FD_1791 port map( D => d(23), CK => n3, RESET => reset, Q => Q(23))
                           ;
   D_I_24 : FD_1790 port map( D => d(24), CK => n3, RESET => reset, Q => Q(24))
                           ;
   D_I_25 : FD_1789 port map( D => d(25), CK => n3, RESET => reset, Q => Q(25))
                           ;
   D_I_26 : FD_1788 port map( D => d(26), CK => n3, RESET => reset, Q => Q(26))
                           ;
   D_I_27 : FD_1787 port map( D => d(27), CK => n3, RESET => reset, Q => Q(27))
                           ;
   D_I_28 : FD_1786 port map( D => d(28), CK => n3, RESET => reset, Q => Q(28))
                           ;
   D_I_29 : FD_1785 port map( D => d(29), CK => n3, RESET => reset, Q => Q(29))
                           ;
   D_I_30 : FD_1784 port map( D => d(30), CK => n3, RESET => reset, Q => Q(30))
                           ;
   D_I_31 : FD_1783 port map( D => d(31), CK => n3, RESET => reset, Q => Q(31))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n1);
   U2 : BUF_X1 port map( A => clk, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_6 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_6;

architecture SYN_struc of reg_nbit_n32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1751
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1752
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1753
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1754
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1755
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1756
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1757
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1758
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1759
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1760
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1761
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1762
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1763
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1764
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1765
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1766
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1767
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1768
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1769
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1770
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1771
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1772
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1773
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1774
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1775
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1776
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1777
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1778
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1779
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1780
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1781
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1782
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1782 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1781 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1780 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1779 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1778 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1777 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1776 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1775 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1774 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1773 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1772 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1771 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1770 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1769 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1768 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1767 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1766 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1765 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1764 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1763 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1762 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1761 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1760 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1759 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1758 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1757 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1756 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1755 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1754 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1753 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1752 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1751 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_5 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_5;

architecture SYN_struc of reg_nbit_n32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1470
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1471
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1472
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1473
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1474
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1475
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1476
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1477
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1478
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1479
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1480
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1481
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1482
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1483
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1484
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1485
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1486
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1487
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1488
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1489
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1490
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1491
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1492
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1493
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1494
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1495
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1496
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1497
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1498
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1499
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1500
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1501
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1501 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1500 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1499 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1498 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1497 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1496 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1495 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1494 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1493 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1492 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1491 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1490 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1489 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1488 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1487 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1486 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1485 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1484 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1483 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1482 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1481 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1480 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1479 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1478 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1477 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1476 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1475 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1474 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1473 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1472 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1471 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1470 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_4 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_4;

architecture SYN_struc of reg_nbit_n32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1189
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1190
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1191
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1192
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1193
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1194
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1195
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1196
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1197
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1198
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1199
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1200
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1201
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1202
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1203
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1204
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1205
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1206
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1207
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1208
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1209
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1210
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1211
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1212
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1213
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1214
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1215
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1216
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1217
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1218
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1219
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1220
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1220 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1219 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1218 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1217 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1216 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1215 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1214 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1213 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1212 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1211 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1210 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1209 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1208 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1207 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1206 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1205 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1204 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1203 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1202 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1201 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1200 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1199 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1198 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1197 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1196 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1195 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1194 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1193 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1192 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1191 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1190 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1189 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_3 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_3;

architecture SYN_struc of reg_nbit_n32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_908
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_909
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_910
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_911
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_912
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_913
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_914
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_915
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_916
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_917
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_918
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_919
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_920
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_921
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_922
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_923
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_924
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_925
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_926
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_927
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_928
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_929
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_930
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_931
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_932
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_933
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_934
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_935
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_936
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_937
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_938
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_939
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_939 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_938 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_937 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_936 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_935 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_934 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_933 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_932 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_931 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_930 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_929 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_928 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_927 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_926 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_925 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_924 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_923 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_922 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_921 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_920 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_919 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_918 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_917 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_916 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_915 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_914 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_913 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_912 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_911 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_910 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_909 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_908 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_2 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_2;

architecture SYN_struc of reg_nbit_n32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_627
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_628
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_629
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_630
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_631
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_632
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_633
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_634
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_635
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_636
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_637
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_638
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_639
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_640
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_641
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_642
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_643
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_644
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_645
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_646
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_647
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_648
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_649
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_650
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_651
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_652
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_653
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_654
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_655
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_656
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_657
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_658
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_658 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_657 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_656 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_655 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_654 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_653 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_652 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_651 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_650 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_649 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_648 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_647 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_646 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_645 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_644 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_643 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_642 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_641 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_640 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_639 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_638 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_637 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_636 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_635 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_634 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_633 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_632 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_631 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_630 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_629 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_628 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_627 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_1;

architecture SYN_struc of reg_nbit_n32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_346
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_347
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_348
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_349
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_350
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_351
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_352
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_353
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_354
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_355
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_356
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_357
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_358
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_359
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_360
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_361
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_362
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_363
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_364
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_365
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_366
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_367
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_368
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_369
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_370
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_371
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_372
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_373
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_374
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_375
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_376
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_377
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_377 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_376 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_375 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_374 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_373 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_372 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_371 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_370 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_369 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_368 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_367 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_366 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_365 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_364 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_363 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_362 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_361 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_360 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_359 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_358 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_357 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_356 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_355 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_354 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_353 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_352 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_351 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_350 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_349 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_348 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_347 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_346 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2249 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2249;

architecture SYN_PLUTO of FD_2249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1098 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1098);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2248 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2248;

architecture SYN_PLUTO of FD_2248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1099 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1099);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2247 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2247;

architecture SYN_PLUTO of FD_2247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1100 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1100);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2246 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2246;

architecture SYN_PLUTO of FD_2246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1101 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1101);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2245 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2245;

architecture SYN_PLUTO of FD_2245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1102 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1102);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2244 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2244;

architecture SYN_PLUTO of FD_2244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1103 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1103);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2243 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2243;

architecture SYN_PLUTO of FD_2243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1104 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1104);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2242 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2242;

architecture SYN_PLUTO of FD_2242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1105 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1105);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2241 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2241;

architecture SYN_PLUTO of FD_2241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1106 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1106);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2240 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2240;

architecture SYN_PLUTO of FD_2240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1107 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1107);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2239 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2239;

architecture SYN_PLUTO of FD_2239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1108 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1108);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2238 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2238;

architecture SYN_PLUTO of FD_2238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1109 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1109);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2237 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2237;

architecture SYN_PLUTO of FD_2237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1110 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1110);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2236 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2236;

architecture SYN_PLUTO of FD_2236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1111 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1111);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2235 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2235;

architecture SYN_PLUTO of FD_2235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1112 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1112);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2234 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2234;

architecture SYN_PLUTO of FD_2234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1113 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1113);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2233 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2233;

architecture SYN_PLUTO of FD_2233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1114 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1114);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2232 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2232;

architecture SYN_PLUTO of FD_2232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1115 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1115);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2231 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2231;

architecture SYN_PLUTO of FD_2231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1116 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1116);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2230 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2230;

architecture SYN_PLUTO of FD_2230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1117 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1117);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2229 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2229;

architecture SYN_PLUTO of FD_2229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1118 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1118);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2228 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2228;

architecture SYN_PLUTO of FD_2228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1119 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1119);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2227 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2227;

architecture SYN_PLUTO of FD_2227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1120 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1120);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2226 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2226;

architecture SYN_PLUTO of FD_2226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1121 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1121);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2225 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2225;

architecture SYN_PLUTO of FD_2225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1122 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1122);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2224 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2224;

architecture SYN_PLUTO of FD_2224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1123 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1123);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2223 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2223;

architecture SYN_PLUTO of FD_2223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1124 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1124);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2222 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2222;

architecture SYN_PLUTO of FD_2222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1125 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1125);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2221 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2221;

architecture SYN_PLUTO of FD_2221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1126 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1126);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2220 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2220;

architecture SYN_PLUTO of FD_2220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1127 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1127);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2219 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2219;

architecture SYN_PLUTO of FD_2219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1128 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1128);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2218 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2218;

architecture SYN_PLUTO of FD_2218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1129 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1129);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2217 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2217;

architecture SYN_PLUTO of FD_2217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1130 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1130);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2216 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2216;

architecture SYN_PLUTO of FD_2216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1131 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1131);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2215 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2215;

architecture SYN_PLUTO of FD_2215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1132 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1132);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2214 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2214;

architecture SYN_PLUTO of FD_2214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1133 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1133);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2213 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2213;

architecture SYN_PLUTO of FD_2213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1134 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1134);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2212 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2212;

architecture SYN_PLUTO of FD_2212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1135 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1135);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2211 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2211;

architecture SYN_PLUTO of FD_2211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1136 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1136);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2210 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2210;

architecture SYN_PLUTO of FD_2210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1137 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1137);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2209 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2209;

architecture SYN_PLUTO of FD_2209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1138 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1138);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2208 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2208;

architecture SYN_PLUTO of FD_2208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1139 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1139);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2207 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2207;

architecture SYN_PLUTO of FD_2207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1140 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1140);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2206 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2206;

architecture SYN_PLUTO of FD_2206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1141 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1141);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2205 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2205;

architecture SYN_PLUTO of FD_2205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1142 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1142);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2204 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2204;

architecture SYN_PLUTO of FD_2204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1143 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1143);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2203 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2203;

architecture SYN_PLUTO of FD_2203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1144 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1144);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2202 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2202;

architecture SYN_PLUTO of FD_2202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1145 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1145);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2201 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2201;

architecture SYN_PLUTO of FD_2201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1146 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1146);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2200 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2200;

architecture SYN_PLUTO of FD_2200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1147 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1147);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2199 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2199;

architecture SYN_PLUTO of FD_2199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1148 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1148);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2198 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2198;

architecture SYN_PLUTO of FD_2198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1149 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1149);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2197 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2197;

architecture SYN_PLUTO of FD_2197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1150 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1150);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2196 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2196;

architecture SYN_PLUTO of FD_2196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1151 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1151);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2195 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2195;

architecture SYN_PLUTO of FD_2195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1152 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1152);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2194 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2194;

architecture SYN_PLUTO of FD_2194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1153 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1153);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2193 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2193;

architecture SYN_PLUTO of FD_2193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1154 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1154);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2192 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2192;

architecture SYN_PLUTO of FD_2192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1155 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1155);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2191 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2191;

architecture SYN_PLUTO of FD_2191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1156 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1156);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2190 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2190;

architecture SYN_PLUTO of FD_2190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1157 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1157);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2189 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2189;

architecture SYN_PLUTO of FD_2189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1158 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1158);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2188 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2188;

architecture SYN_PLUTO of FD_2188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1159 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1159);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2187 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2187;

architecture SYN_PLUTO of FD_2187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1160 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1160);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2186 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2186;

architecture SYN_PLUTO of FD_2186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1161 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1161);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2185 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2185;

architecture SYN_PLUTO of FD_2185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1162 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1162);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2184 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2184;

architecture SYN_PLUTO of FD_2184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1163 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1163);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2183 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2183;

architecture SYN_PLUTO of FD_2183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1164 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1164);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2182 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2182;

architecture SYN_PLUTO of FD_2182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1165 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1165);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2181 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2181;

architecture SYN_PLUTO of FD_2181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1166 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1166);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2180 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2180;

architecture SYN_PLUTO of FD_2180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1167 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1167);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2179 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2179;

architecture SYN_PLUTO of FD_2179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1168 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1168);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2178 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2178;

architecture SYN_PLUTO of FD_2178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1169 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1169);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2177 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2177;

architecture SYN_PLUTO of FD_2177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1170 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1170);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2176 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2176;

architecture SYN_PLUTO of FD_2176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1171 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1171);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2175 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2175;

architecture SYN_PLUTO of FD_2175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1172 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1172);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2174 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2174;

architecture SYN_PLUTO of FD_2174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1173 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1173);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2173 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2173;

architecture SYN_PLUTO of FD_2173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1174 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1174);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2172 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2172;

architecture SYN_PLUTO of FD_2172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1175 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1175);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2171 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2171;

architecture SYN_PLUTO of FD_2171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1176 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1176);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2170 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2170;

architecture SYN_PLUTO of FD_2170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1177 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1177);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2169 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2169;

architecture SYN_PLUTO of FD_2169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1178 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1178);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2168 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2168;

architecture SYN_PLUTO of FD_2168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1179 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1179);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2167 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2167;

architecture SYN_PLUTO of FD_2167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1180 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1180);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2166 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2166;

architecture SYN_PLUTO of FD_2166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1181 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1181);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2165 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2165;

architecture SYN_PLUTO of FD_2165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1182 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1182);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2164 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2164;

architecture SYN_PLUTO of FD_2164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1183 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1183);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2163 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2163;

architecture SYN_PLUTO of FD_2163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1184 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1184);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2162 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2162;

architecture SYN_PLUTO of FD_2162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1185 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1185);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2161 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2161;

architecture SYN_PLUTO of FD_2161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1186 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1186);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2160 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2160;

architecture SYN_PLUTO of FD_2160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1187 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1187);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2159 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2159;

architecture SYN_PLUTO of FD_2159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1188 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1188);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2158 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2158;

architecture SYN_PLUTO of FD_2158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1189 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1189);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2157 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2157;

architecture SYN_PLUTO of FD_2157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1190 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1190);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2156 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2156;

architecture SYN_PLUTO of FD_2156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1191 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1191);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2155 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2155;

architecture SYN_PLUTO of FD_2155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1192 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1192);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2154 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2154;

architecture SYN_PLUTO of FD_2154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1193 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1193);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2153 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2153;

architecture SYN_PLUTO of FD_2153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1194 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1194);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2152 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2152;

architecture SYN_PLUTO of FD_2152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1195 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1195);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2151 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2151;

architecture SYN_PLUTO_architecture of FD_2151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1196 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1196);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2150 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2150;

architecture SYN_PLUTO_architecture2 of FD_2150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1197 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1197);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2149 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2149;

architecture SYN_PLUTO_architecture3 of FD_2149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1198 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1198);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2148 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2148;

architecture SYN_PLUTO_architecture4 of FD_2148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1199 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1199);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2147 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2147;

architecture SYN_PLUTO_architecture5 of FD_2147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1200 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1200);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2146 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2146;

architecture SYN_PLUTO_architecture6 of FD_2146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1201 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1201);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2145 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2145;

architecture SYN_PLUTO_architecture7 of FD_2145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1202 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1202);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2144 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2144;

architecture SYN_PLUTO_architecture8 of FD_2144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1203 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1203);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2143 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2143;

architecture SYN_PLUTO_architecture9 of FD_2143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1204 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1204);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2142 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2142;

architecture SYN_PLUTO_architecture10 of FD_2142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1205 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1205);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2141 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2141;

architecture SYN_PLUTO_architecture11 of FD_2141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1206 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1206);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2140 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2140;

architecture SYN_PLUTO_architecture12 of FD_2140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1207 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1207);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2139 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2139;

architecture SYN_PLUTO_architecture13 of FD_2139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1208 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1208);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2138 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2138;

architecture SYN_PLUTO_architecture14 of FD_2138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1209 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1209);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2137 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2137;

architecture SYN_PLUTO_architecture15 of FD_2137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1210 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1210);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2136 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2136;

architecture SYN_PLUTO_architecture16 of FD_2136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1211 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1211);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2135 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2135;

architecture SYN_PLUTO_architecture17 of FD_2135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1212 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1212);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2134 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2134;

architecture SYN_PLUTO_architecture18 of FD_2134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1213 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1213);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2133 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2133;

architecture SYN_PLUTO_architecture19 of FD_2133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1214 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1214);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2132 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2132;

architecture SYN_PLUTO_architecture20 of FD_2132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1215 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1215);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2131 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2131;

architecture SYN_PLUTO_architecture21 of FD_2131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1216 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1216);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2130 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2130;

architecture SYN_PLUTO_architecture22 of FD_2130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1217 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1217);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2129 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2129;

architecture SYN_PLUTO_architecture23 of FD_2129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1218 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1218);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2128 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2128;

architecture SYN_PLUTO_architecture24 of FD_2128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1219 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1219);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2127 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2127;

architecture SYN_PLUTO_architecture25 of FD_2127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1220 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1220);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2126 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2126;

architecture SYN_PLUTO_architecture26 of FD_2126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1221 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1221);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2125 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2125;

architecture SYN_PLUTO_architecture27 of FD_2125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1222 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1222);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2124 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2124;

architecture SYN_PLUTO_architecture28 of FD_2124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1223 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1223);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2123 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2123;

architecture SYN_PLUTO_architecture29 of FD_2123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1224 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1224);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2122 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2122;

architecture SYN_PLUTO_architecture30 of FD_2122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1225 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1225);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2121 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2121;

architecture SYN_PLUTO_architecture31 of FD_2121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1226 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1226);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2120 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2120;

architecture SYN_PLUTO of FD_2120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1227 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1227);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2119 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2119;

architecture SYN_PLUTO_architecture of FD_2119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1228 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1228);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2118 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2118;

architecture SYN_PLUTO_architecture2 of FD_2118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1229 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1229);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2117 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2117;

architecture SYN_PLUTO_architecture3 of FD_2117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1230 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1230);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2116 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2116;

architecture SYN_PLUTO_architecture4 of FD_2116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1231 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1231);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2115 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2115;

architecture SYN_PLUTO_architecture5 of FD_2115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1232 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1232);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2114 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2114;

architecture SYN_PLUTO_architecture6 of FD_2114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1233 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1233);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2113 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2113;

architecture SYN_PLUTO_architecture7 of FD_2113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1234 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1234);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2112 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2112;

architecture SYN_PLUTO_architecture8 of FD_2112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1235 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1235);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2111 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2111;

architecture SYN_PLUTO_architecture9 of FD_2111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1236 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1236);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2110 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2110;

architecture SYN_PLUTO_architecture10 of FD_2110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1237 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1237);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2109 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2109;

architecture SYN_PLUTO_architecture11 of FD_2109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1238 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1238);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2108 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2108;

architecture SYN_PLUTO_architecture12 of FD_2108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1239 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1239);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2107 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2107;

architecture SYN_PLUTO_architecture13 of FD_2107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1240 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1240);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2106 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2106;

architecture SYN_PLUTO_architecture14 of FD_2106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1241 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1241);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2105 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2105;

architecture SYN_PLUTO_architecture15 of FD_2105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1242 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1242);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2104 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2104;

architecture SYN_PLUTO_architecture16 of FD_2104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1243 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1243);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2103 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2103;

architecture SYN_PLUTO_architecture17 of FD_2103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1244 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1244);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2102 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2102;

architecture SYN_PLUTO_architecture18 of FD_2102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1245 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1245);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2101 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2101;

architecture SYN_PLUTO_architecture19 of FD_2101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1246 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1246);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2100 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2100;

architecture SYN_PLUTO_architecture20 of FD_2100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1247 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1247);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2099 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2099;

architecture SYN_PLUTO_architecture21 of FD_2099 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1248 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1248);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2098 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2098;

architecture SYN_PLUTO_architecture22 of FD_2098 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1249 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1249);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2097 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2097;

architecture SYN_PLUTO_architecture23 of FD_2097 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1250 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1250);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2096 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2096;

architecture SYN_PLUTO_architecture24 of FD_2096 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1251 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1251);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2095 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2095;

architecture SYN_PLUTO_architecture25 of FD_2095 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1252 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1252);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2094 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2094;

architecture SYN_PLUTO_architecture26 of FD_2094 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1253 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1253);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2093 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2093;

architecture SYN_PLUTO_architecture27 of FD_2093 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1254 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1254);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2092 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2092;

architecture SYN_PLUTO_architecture28 of FD_2092 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1255 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1255);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2091 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2091;

architecture SYN_PLUTO_architecture29 of FD_2091 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1256 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1256);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2090 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2090;

architecture SYN_PLUTO_architecture30 of FD_2090 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1257 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1257);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2089 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2089;

architecture SYN_PLUTO_architecture31 of FD_2089 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1258 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1258);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2088 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2088;

architecture SYN_PLUTO of FD_2088 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1259 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1259);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2087 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2087;

architecture SYN_PLUTO of FD_2087 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1260 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1260);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2086 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2086;

architecture SYN_PLUTO of FD_2086 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1261 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1261);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2085 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2085;

architecture SYN_PLUTO of FD_2085 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1262 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1262);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2084 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2084;

architecture SYN_PLUTO of FD_2084 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1263 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1263);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2083 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2083;

architecture SYN_PLUTO of FD_2083 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1264 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1264);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2082 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2082;

architecture SYN_PLUTO_architecture of FD_2082 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1265 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1265);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2081 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2081;

architecture SYN_PLUTO_architecture2 of FD_2081 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1266 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1266);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2080 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2080;

architecture SYN_PLUTO_architecture3 of FD_2080 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1267 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1267);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2079 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2079;

architecture SYN_PLUTO_architecture4 of FD_2079 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1268 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1268);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2078 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2078;

architecture SYN_PLUTO of FD_2078 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1269 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1269);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2077 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2077;

architecture SYN_PLUTO_architecture of FD_2077 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1270 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1270);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2076 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2076;

architecture SYN_PLUTO_architecture2 of FD_2076 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1271 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1271);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2075 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2075;

architecture SYN_PLUTO_architecture3 of FD_2075 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1272 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1272);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2074 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2074;

architecture SYN_PLUTO_architecture4 of FD_2074 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1273 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1273);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2073 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2073;

architecture SYN_PLUTO of FD_2073 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1274 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1274);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2072 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2072;

architecture SYN_PLUTO_architecture of FD_2072 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1275 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1275);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2071 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2071;

architecture SYN_PLUTO_architecture2 of FD_2071 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1276 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1276);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2070 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2070;

architecture SYN_PLUTO_architecture3 of FD_2070 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1277 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1277);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2069 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2069;

architecture SYN_PLUTO_architecture4 of FD_2069 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1278 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1278);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2068 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2068;

architecture SYN_PLUTO_architecture5 of FD_2068 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1279 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1279);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2067 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2067;

architecture SYN_PLUTO_architecture6 of FD_2067 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1280 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1280);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2066 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2066;

architecture SYN_PLUTO_architecture7 of FD_2066 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1281 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1281);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2065 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2065;

architecture SYN_PLUTO_architecture8 of FD_2065 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1282 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1282);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2064 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2064;

architecture SYN_PLUTO_architecture9 of FD_2064 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1283 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1283);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2063 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2063;

architecture SYN_PLUTO_architecture10 of FD_2063 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1284 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1284);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2062 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2062;

architecture SYN_PLUTO_architecture11 of FD_2062 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1285 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1285);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2061 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2061;

architecture SYN_PLUTO_architecture12 of FD_2061 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1286 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1286);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2060 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2060;

architecture SYN_PLUTO_architecture13 of FD_2060 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1287 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1287);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2059 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2059;

architecture SYN_PLUTO_architecture14 of FD_2059 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1288 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1288);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2058 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2058;

architecture SYN_PLUTO_architecture15 of FD_2058 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1289 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1289);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2057 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2057;

architecture SYN_PLUTO_architecture16 of FD_2057 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1290 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1290);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2056 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2056;

architecture SYN_PLUTO_architecture17 of FD_2056 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1291 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1291);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2055 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2055;

architecture SYN_PLUTO_architecture18 of FD_2055 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1292 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1292);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2054 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2054;

architecture SYN_PLUTO_architecture19 of FD_2054 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1293 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1293);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2053 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2053;

architecture SYN_PLUTO_architecture20 of FD_2053 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1294 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1294);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2052 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2052;

architecture SYN_PLUTO_architecture21 of FD_2052 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1295 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1295);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2051 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2051;

architecture SYN_PLUTO_architecture22 of FD_2051 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1296 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1296);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2050 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2050;

architecture SYN_PLUTO_architecture23 of FD_2050 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1297 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1297);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2049 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2049;

architecture SYN_PLUTO_architecture24 of FD_2049 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1298 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1298);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2048 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2048;

architecture SYN_PLUTO_architecture25 of FD_2048 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1299 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1299);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2047 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2047;

architecture SYN_PLUTO_architecture26 of FD_2047 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1300 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1300);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2046 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2046;

architecture SYN_PLUTO_architecture27 of FD_2046 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1301 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1301);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2045 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2045;

architecture SYN_PLUTO_architecture28 of FD_2045 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1302 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1302);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2044 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2044;

architecture SYN_PLUTO_architecture29 of FD_2044 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1303 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1303);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2043 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2043;

architecture SYN_PLUTO_architecture30 of FD_2043 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1304 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1304);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2042 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2042;

architecture SYN_PLUTO_architecture31 of FD_2042 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1305 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1305);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2041 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2041;

architecture SYN_PLUTO of FD_2041 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1306 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1306);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2040 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2040;

architecture SYN_PLUTO_architecture of FD_2040 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1307 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1307);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2039 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2039;

architecture SYN_PLUTO_architecture2 of FD_2039 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1308 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1308);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2038 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2038;

architecture SYN_PLUTO_architecture3 of FD_2038 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1309 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1309);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2037 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2037;

architecture SYN_PLUTO_architecture4 of FD_2037 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1310 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1310);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2036 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2036;

architecture SYN_PLUTO_architecture5 of FD_2036 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1311 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1311);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2035 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2035;

architecture SYN_PLUTO_architecture6 of FD_2035 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1312 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1312);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2034 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2034;

architecture SYN_PLUTO_architecture7 of FD_2034 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1313 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1313);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2033 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2033;

architecture SYN_PLUTO_architecture8 of FD_2033 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1314 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1314);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2032 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2032;

architecture SYN_PLUTO_architecture9 of FD_2032 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1315 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1315);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2031 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2031;

architecture SYN_PLUTO_architecture10 of FD_2031 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1316 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1316);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2030 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2030;

architecture SYN_PLUTO_architecture11 of FD_2030 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1317 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1317);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2029 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2029;

architecture SYN_PLUTO_architecture12 of FD_2029 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1318 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1318);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2028 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2028;

architecture SYN_PLUTO_architecture13 of FD_2028 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1319 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1319);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2027 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2027;

architecture SYN_PLUTO_architecture14 of FD_2027 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1320 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1320);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2026 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2026;

architecture SYN_PLUTO_architecture15 of FD_2026 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1321 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1321);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2025 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2025;

architecture SYN_PLUTO_architecture16 of FD_2025 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1322 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1322);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2024 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2024;

architecture SYN_PLUTO_architecture17 of FD_2024 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1323 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1323);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2023 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2023;

architecture SYN_PLUTO_architecture18 of FD_2023 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1324 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1324);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2022 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2022;

architecture SYN_PLUTO_architecture19 of FD_2022 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1325 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1325);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2021 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2021;

architecture SYN_PLUTO_architecture20 of FD_2021 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1326 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1326);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2020 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2020;

architecture SYN_PLUTO_architecture21 of FD_2020 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1327 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1327);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2019 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2019;

architecture SYN_PLUTO_architecture22 of FD_2019 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1328 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1328);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2018 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2018;

architecture SYN_PLUTO_architecture23 of FD_2018 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1329 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1329);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2017 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2017;

architecture SYN_PLUTO_architecture24 of FD_2017 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1330 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1330);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2016 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2016;

architecture SYN_PLUTO_architecture25 of FD_2016 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1331 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1331);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2015 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2015;

architecture SYN_PLUTO_architecture26 of FD_2015 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1332 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1332);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2014 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2014;

architecture SYN_PLUTO_architecture27 of FD_2014 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1333 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1333);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2013 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2013;

architecture SYN_PLUTO_architecture28 of FD_2013 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1334 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1334);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2012 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2012;

architecture SYN_PLUTO_architecture29 of FD_2012 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1335 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1335);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2011 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2011;

architecture SYN_PLUTO_architecture30 of FD_2011 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1336 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1336);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2010 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2010;

architecture SYN_PLUTO_architecture31 of FD_2010 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1337 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1337);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2009 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2009;

architecture SYN_PLUTO of FD_2009 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1338 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1338);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2008 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2008;

architecture SYN_PLUTO_architecture of FD_2008 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1339 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1339);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2007 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2007;

architecture SYN_PLUTO_architecture2 of FD_2007 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1340 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1340);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2006 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2006;

architecture SYN_PLUTO_architecture3 of FD_2006 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1341 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1341);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2005 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2005;

architecture SYN_PLUTO_architecture4 of FD_2005 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1342 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1342);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2004 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2004;

architecture SYN_PLUTO_architecture5 of FD_2004 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1343 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1343);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2003 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2003;

architecture SYN_PLUTO_architecture6 of FD_2003 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1344 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1344);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2002 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2002;

architecture SYN_PLUTO_architecture7 of FD_2002 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1345 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1345);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2001 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2001;

architecture SYN_PLUTO_architecture8 of FD_2001 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1346 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1346);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2000 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2000;

architecture SYN_PLUTO_architecture9 of FD_2000 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1347 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1347);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1999 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1999;

architecture SYN_PLUTO_architecture10 of FD_1999 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1348 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1348);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1998 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1998;

architecture SYN_PLUTO_architecture11 of FD_1998 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1349 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1349);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1997 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1997;

architecture SYN_PLUTO_architecture12 of FD_1997 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1350 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1350);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1996 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1996;

architecture SYN_PLUTO_architecture13 of FD_1996 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1351 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1351);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1995 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1995;

architecture SYN_PLUTO_architecture14 of FD_1995 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1352 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1352);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1994 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1994;

architecture SYN_PLUTO_architecture15 of FD_1994 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1353 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1353);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1993 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1993;

architecture SYN_PLUTO_architecture16 of FD_1993 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1354 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1354);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1992 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1992;

architecture SYN_PLUTO_architecture17 of FD_1992 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1355 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1355);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1991 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1991;

architecture SYN_PLUTO_architecture18 of FD_1991 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1356 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1356);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1990 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1990;

architecture SYN_PLUTO_architecture19 of FD_1990 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1357 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1357);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1989 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1989;

architecture SYN_PLUTO_architecture20 of FD_1989 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1358 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1358);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1988 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1988;

architecture SYN_PLUTO_architecture21 of FD_1988 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1359 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1359);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1987 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1987;

architecture SYN_PLUTO_architecture22 of FD_1987 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1360 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1360);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1986 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1986;

architecture SYN_PLUTO_architecture23 of FD_1986 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1361 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1361);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1985 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1985;

architecture SYN_PLUTO_architecture24 of FD_1985 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1362 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1362);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1984 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1984;

architecture SYN_PLUTO_architecture25 of FD_1984 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1363 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1363);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1983 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1983;

architecture SYN_PLUTO_architecture26 of FD_1983 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1364 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1364);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1982 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1982;

architecture SYN_PLUTO_architecture27 of FD_1982 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1365 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1365);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1981 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1981;

architecture SYN_PLUTO_architecture28 of FD_1981 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1366 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1366);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1980 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1980;

architecture SYN_PLUTO_architecture29 of FD_1980 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1367 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1367);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1979 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1979;

architecture SYN_PLUTO_architecture30 of FD_1979 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1368 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1368);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1978 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1978;

architecture SYN_PLUTO_architecture31 of FD_1978 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1369 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1369);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1977 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1977;

architecture SYN_PLUTO of FD_1977 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1370 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1370);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1976 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1976;

architecture SYN_PLUTO of FD_1976 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1371 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1371);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1975 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1975;

architecture SYN_PLUTO of FD_1975 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1372 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1372);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1974 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1974;

architecture SYN_PLUTO of FD_1974 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1373 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1373);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1973 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1973;

architecture SYN_PLUTO of FD_1973 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1374 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1374);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1972 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1972;

architecture SYN_PLUTO of FD_1972 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1375 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1375);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1971 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1971;

architecture SYN_PLUTO of FD_1971 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1376 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1376);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1970 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1970;

architecture SYN_PLUTO of FD_1970 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1377 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1377);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1969 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1969;

architecture SYN_PLUTO of FD_1969 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1378 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1378);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1968 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1968;

architecture SYN_PLUTO of FD_1968 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1379 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1379);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1967 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1967;

architecture SYN_PLUTO of FD_1967 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1380 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1380);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1966 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1966;

architecture SYN_PLUTO of FD_1966 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1381 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1381);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1965 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1965;

architecture SYN_PLUTO of FD_1965 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1382 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1382);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1964 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1964;

architecture SYN_PLUTO of FD_1964 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1383 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1383);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1963 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1963;

architecture SYN_PLUTO of FD_1963 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1384 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1384);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1962 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1962;

architecture SYN_PLUTO of FD_1962 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1385 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1385);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1961 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1961;

architecture SYN_PLUTO of FD_1961 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1386 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1386);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1960 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1960;

architecture SYN_PLUTO of FD_1960 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1387 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1387);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1959 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1959;

architecture SYN_PLUTO of FD_1959 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1388 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1388);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1958 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1958;

architecture SYN_PLUTO of FD_1958 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1389 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1389);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1957 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1957;

architecture SYN_PLUTO of FD_1957 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1390 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1390);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1956 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1956;

architecture SYN_PLUTO of FD_1956 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1391 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1391);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1955 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1955;

architecture SYN_PLUTO of FD_1955 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1392 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1392);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1954 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1954;

architecture SYN_PLUTO of FD_1954 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1393 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1393);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1953 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1953;

architecture SYN_PLUTO of FD_1953 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1394 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1394);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1952 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1952;

architecture SYN_PLUTO of FD_1952 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1395 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1395);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1951 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1951;

architecture SYN_PLUTO of FD_1951 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1396 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1396);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1950 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1950;

architecture SYN_PLUTO of FD_1950 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1397 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1397);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1949 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1949;

architecture SYN_PLUTO of FD_1949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1398 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1398);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1948 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1948;

architecture SYN_PLUTO of FD_1948 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1399 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1399);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1947 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1947;

architecture SYN_PLUTO of FD_1947 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1400 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1400);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1946 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1946;

architecture SYN_PLUTO of FD_1946 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1401 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1401);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1945 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1945;

architecture SYN_PLUTO of FD_1945 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1402 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1402);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1944 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1944;

architecture SYN_PLUTO of FD_1944 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1403 : std_logic;

begin
   
   Q_reg : DFFR_X2 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1403);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1943 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1943;

architecture SYN_PLUTO_architecture of FD_1943 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1404 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1404);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1942 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1942;

architecture SYN_PLUTO_architecture2 of FD_1942 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1405 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1405);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1941 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1941;

architecture SYN_PLUTO_architecture3 of FD_1941 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1406 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1406);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1940 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1940;

architecture SYN_PLUTO_architecture4 of FD_1940 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1407 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1407);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1939 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1939;

architecture SYN_PLUTO_architecture5 of FD_1939 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1408 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1408);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1938 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1938;

architecture SYN_PLUTO_architecture6 of FD_1938 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1409 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1409);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1937 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1937;

architecture SYN_PLUTO_architecture7 of FD_1937 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1410 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1410);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1936 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1936;

architecture SYN_PLUTO_architecture8 of FD_1936 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1411 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1411);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1935 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1935;

architecture SYN_PLUTO_architecture9 of FD_1935 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1412 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1412);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1934 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1934;

architecture SYN_PLUTO_architecture10 of FD_1934 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1413 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1413);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1933 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1933;

architecture SYN_PLUTO_architecture11 of FD_1933 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1414 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1414);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1932 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1932;

architecture SYN_PLUTO_architecture12 of FD_1932 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1415 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1415);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1931 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1931;

architecture SYN_PLUTO_architecture13 of FD_1931 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1416 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1416);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1930 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1930;

architecture SYN_PLUTO_architecture14 of FD_1930 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1417 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1417);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1929 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1929;

architecture SYN_PLUTO_architecture15 of FD_1929 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1418 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1418);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1928 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1928;

architecture SYN_PLUTO_architecture16 of FD_1928 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1419 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1419);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1927 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1927;

architecture SYN_PLUTO_architecture17 of FD_1927 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1420 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1420);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1926 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1926;

architecture SYN_PLUTO_architecture18 of FD_1926 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1421 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1421);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1925 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1925;

architecture SYN_PLUTO_architecture19 of FD_1925 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1422 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1422);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1924 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1924;

architecture SYN_PLUTO_architecture20 of FD_1924 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1423 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1423);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1923 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1923;

architecture SYN_PLUTO_architecture21 of FD_1923 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1424 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1424);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1922 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1922;

architecture SYN_PLUTO_architecture22 of FD_1922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1425 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1425);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1921 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1921;

architecture SYN_PLUTO_architecture23 of FD_1921 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1426 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1426);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1920 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1920;

architecture SYN_PLUTO_architecture24 of FD_1920 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1427 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1427);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1919 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1919;

architecture SYN_PLUTO_architecture25 of FD_1919 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1428 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1428);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1918 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1918;

architecture SYN_PLUTO_architecture26 of FD_1918 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1429 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1429);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1917 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1917;

architecture SYN_PLUTO_architecture27 of FD_1917 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1430 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1430);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1916 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1916;

architecture SYN_PLUTO_architecture28 of FD_1916 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1431 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1431);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1915 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1915;

architecture SYN_PLUTO_architecture29 of FD_1915 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1432 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1432);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1914 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1914;

architecture SYN_PLUTO_architecture30 of FD_1914 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1433 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1433);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1913 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1913;

architecture SYN_PLUTO_architecture31 of FD_1913 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1434 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1434);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1912 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1912;

architecture SYN_PLUTO_architecture32 of FD_1912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1435 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1435);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1911 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1911;

architecture SYN_PLUTO of FD_1911 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1436 : std_logic;

begin
   
   Q_reg : DFFR_X2 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1436);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1910 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1910;

architecture SYN_PLUTO of FD_1910 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1437 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1437);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1909 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1909;

architecture SYN_PLUTO_architecture of FD_1909 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1438 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1438);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1908 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1908;

architecture SYN_PLUTO_architecture2 of FD_1908 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1439 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1439);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1907 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1907;

architecture SYN_PLUTO_architecture3 of FD_1907 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1440 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1440);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1906 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1906;

architecture SYN_PLUTO_architecture4 of FD_1906 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1441 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1441);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1905 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1905;

architecture SYN_PLUTO_architecture5 of FD_1905 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1442 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1442);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1904 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1904;

architecture SYN_PLUTO_architecture6 of FD_1904 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1443 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1443);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1903 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1903;

architecture SYN_PLUTO_architecture7 of FD_1903 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1444 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1444);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1902 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1902;

architecture SYN_PLUTO_architecture8 of FD_1902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1445 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1445);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1901 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1901;

architecture SYN_PLUTO_architecture9 of FD_1901 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1446 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1446);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1900 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1900;

architecture SYN_PLUTO_architecture10 of FD_1900 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1447 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1447);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1899 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1899;

architecture SYN_PLUTO_architecture11 of FD_1899 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1448 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1448);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1898 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1898;

architecture SYN_PLUTO_architecture12 of FD_1898 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1449 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1449);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1897 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1897;

architecture SYN_PLUTO_architecture13 of FD_1897 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1450 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1450);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1896 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1896;

architecture SYN_PLUTO_architecture14 of FD_1896 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1451 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1451);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1895 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1895;

architecture SYN_PLUTO_architecture15 of FD_1895 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1452 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1452);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1894 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1894;

architecture SYN_PLUTO_architecture16 of FD_1894 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1453 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1453);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1893 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1893;

architecture SYN_PLUTO_architecture17 of FD_1893 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1454 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1454);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1892 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1892;

architecture SYN_PLUTO_architecture18 of FD_1892 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1455 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1455);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1891 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1891;

architecture SYN_PLUTO_architecture19 of FD_1891 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1456 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1456);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1890 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1890;

architecture SYN_PLUTO_architecture20 of FD_1890 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1457 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1457);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1889 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1889;

architecture SYN_PLUTO_architecture21 of FD_1889 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1458 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1458);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1888 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1888;

architecture SYN_PLUTO_architecture22 of FD_1888 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1459 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1459);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1887 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1887;

architecture SYN_PLUTO_architecture23 of FD_1887 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1460 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1460);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1886 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1886;

architecture SYN_PLUTO_architecture24 of FD_1886 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1461 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1461);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1885 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1885;

architecture SYN_PLUTO_architecture25 of FD_1885 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1462 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1462);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1884 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1884;

architecture SYN_PLUTO_architecture26 of FD_1884 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1463 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1463);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1883 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1883;

architecture SYN_PLUTO_architecture27 of FD_1883 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1464 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1464);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1882 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1882;

architecture SYN_PLUTO_architecture28 of FD_1882 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1465 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1465);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1881 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1881;

architecture SYN_PLUTO_architecture29 of FD_1881 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1466 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1466);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1880 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1880;

architecture SYN_PLUTO_architecture30 of FD_1880 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1467 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1467);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1879 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1879;

architecture SYN_PLUTO_architecture31 of FD_1879 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1468 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1468);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1878 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1878;

architecture SYN_PLUTO of FD_1878 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1469 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1469);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1877 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1877;

architecture SYN_PLUTO_architecture of FD_1877 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1470 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1470);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1876 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1876;

architecture SYN_PLUTO_architecture2 of FD_1876 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1471 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1471);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1875 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1875;

architecture SYN_PLUTO_architecture3 of FD_1875 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1472 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1472);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1874 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1874;

architecture SYN_PLUTO_architecture4 of FD_1874 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1473 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1473);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1873 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1873;

architecture SYN_PLUTO_architecture5 of FD_1873 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1474 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1474);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1872 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1872;

architecture SYN_PLUTO_architecture6 of FD_1872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1475 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1475);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1871 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1871;

architecture SYN_PLUTO_architecture7 of FD_1871 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1476 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1476);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1870 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1870;

architecture SYN_PLUTO_architecture8 of FD_1870 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1477 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1477);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1869 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1869;

architecture SYN_PLUTO_architecture9 of FD_1869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1478 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1478);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1868 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1868;

architecture SYN_PLUTO_architecture10 of FD_1868 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1479 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1479);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1867 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1867;

architecture SYN_PLUTO_architecture11 of FD_1867 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1480 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1480);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1866 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1866;

architecture SYN_PLUTO_architecture12 of FD_1866 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1481 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1481);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1865 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1865;

architecture SYN_PLUTO_architecture13 of FD_1865 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1482 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1482);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1864 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1864;

architecture SYN_PLUTO_architecture14 of FD_1864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1483 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1483);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1863 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1863;

architecture SYN_PLUTO_architecture15 of FD_1863 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1484 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1484);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1862 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1862;

architecture SYN_PLUTO_architecture16 of FD_1862 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1485 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1485);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1861 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1861;

architecture SYN_PLUTO_architecture17 of FD_1861 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1486 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1486);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1860 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1860;

architecture SYN_PLUTO_architecture18 of FD_1860 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1487 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1487);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1859 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1859;

architecture SYN_PLUTO_architecture19 of FD_1859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1488 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1488);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1858 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1858;

architecture SYN_PLUTO_architecture20 of FD_1858 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1489 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1489);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1857 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1857;

architecture SYN_PLUTO_architecture21 of FD_1857 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1490 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1490);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1856 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1856;

architecture SYN_PLUTO_architecture22 of FD_1856 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1491 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1491);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1855 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1855;

architecture SYN_PLUTO_architecture23 of FD_1855 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1492 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1492);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1854 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1854;

architecture SYN_PLUTO_architecture24 of FD_1854 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1493 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1493);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1853 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1853;

architecture SYN_PLUTO_architecture25 of FD_1853 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1494 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1494);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1852 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1852;

architecture SYN_PLUTO_architecture26 of FD_1852 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1495 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1495);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1851 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1851;

architecture SYN_PLUTO_architecture27 of FD_1851 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1496 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1496);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1850 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1850;

architecture SYN_PLUTO_architecture28 of FD_1850 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1497 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1497);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1849 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1849;

architecture SYN_PLUTO_architecture29 of FD_1849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1498 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1498);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1848 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1848;

architecture SYN_PLUTO_architecture30 of FD_1848 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1499 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1499);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1847 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1847;

architecture SYN_PLUTO_architecture31 of FD_1847 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1500 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1500);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1846 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1846;

architecture SYN_PLUTO of FD_1846 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1501 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1501);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1845 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1845;

architecture SYN_PLUTO_architecture of FD_1845 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1502 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1502);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1844 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1844;

architecture SYN_PLUTO_architecture2 of FD_1844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1503 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1503);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1843 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1843;

architecture SYN_PLUTO_architecture3 of FD_1843 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1504 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1504);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1842 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1842;

architecture SYN_PLUTO_architecture4 of FD_1842 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1505 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1505);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1841 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1841;

architecture SYN_PLUTO_architecture5 of FD_1841 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1506 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1506);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1840 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1840;

architecture SYN_PLUTO_architecture6 of FD_1840 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1507 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1507);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1839 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1839;

architecture SYN_PLUTO_architecture7 of FD_1839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1508 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1508);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1838 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1838;

architecture SYN_PLUTO_architecture8 of FD_1838 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1509 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1509);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1837 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1837;

architecture SYN_PLUTO_architecture9 of FD_1837 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1510 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1510);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1836 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1836;

architecture SYN_PLUTO_architecture10 of FD_1836 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1511 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1511);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1835 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1835;

architecture SYN_PLUTO_architecture11 of FD_1835 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1512 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1512);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1834 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1834;

architecture SYN_PLUTO_architecture12 of FD_1834 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1513 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1513);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1833 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1833;

architecture SYN_PLUTO_architecture13 of FD_1833 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1514 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1514);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1832 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1832;

architecture SYN_PLUTO_architecture14 of FD_1832 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1515 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1515);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1831 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1831;

architecture SYN_PLUTO_architecture15 of FD_1831 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1516 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1516);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1830 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1830;

architecture SYN_PLUTO_architecture16 of FD_1830 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1517 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1517);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1829 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1829;

architecture SYN_PLUTO_architecture17 of FD_1829 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1518 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1518);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1828 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1828;

architecture SYN_PLUTO_architecture18 of FD_1828 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1519 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1519);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1827 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1827;

architecture SYN_PLUTO_architecture19 of FD_1827 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1520 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1520);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1826 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1826;

architecture SYN_PLUTO_architecture20 of FD_1826 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1521 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1521);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1825 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1825;

architecture SYN_PLUTO_architecture21 of FD_1825 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1522 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1522);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1824 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1824;

architecture SYN_PLUTO_architecture22 of FD_1824 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1523 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1523);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1823 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1823;

architecture SYN_PLUTO_architecture23 of FD_1823 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1524 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1524);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1822 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1822;

architecture SYN_PLUTO_architecture24 of FD_1822 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1525 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1525);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1821 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1821;

architecture SYN_PLUTO_architecture25 of FD_1821 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1526 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1526);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1820 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1820;

architecture SYN_PLUTO_architecture26 of FD_1820 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1527 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1527);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1819 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1819;

architecture SYN_PLUTO_architecture27 of FD_1819 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1528 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1528);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1818 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1818;

architecture SYN_PLUTO_architecture28 of FD_1818 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1529 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1529);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1817 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1817;

architecture SYN_PLUTO_architecture29 of FD_1817 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1530 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1530);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1816 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1816;

architecture SYN_PLUTO_architecture30 of FD_1816 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1531 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1531);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1815 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1815;

architecture SYN_PLUTO_architecture31 of FD_1815 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1532 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1532);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1814 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1814;

architecture SYN_PLUTO of FD_1814 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1533 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1533);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1813 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1813;

architecture SYN_PLUTO_architecture of FD_1813 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1534 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1534);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1812 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1812;

architecture SYN_PLUTO_architecture2 of FD_1812 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1535 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1535);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1811 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1811;

architecture SYN_PLUTO_architecture3 of FD_1811 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1536 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1536);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1810 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1810;

architecture SYN_PLUTO_architecture4 of FD_1810 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1537 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1537);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1809 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1809;

architecture SYN_PLUTO_architecture5 of FD_1809 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1538 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1538);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1808 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1808;

architecture SYN_PLUTO_architecture6 of FD_1808 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1539 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1539);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1807 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1807;

architecture SYN_PLUTO_architecture7 of FD_1807 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1540 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1540);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1806 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1806;

architecture SYN_PLUTO_architecture8 of FD_1806 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1541 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1541);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1805 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1805;

architecture SYN_PLUTO_architecture9 of FD_1805 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1542 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1542);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1804 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1804;

architecture SYN_PLUTO_architecture10 of FD_1804 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1543 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1543);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1803 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1803;

architecture SYN_PLUTO_architecture11 of FD_1803 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1544 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1544);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1802 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1802;

architecture SYN_PLUTO_architecture12 of FD_1802 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1545 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1545);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1801 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1801;

architecture SYN_PLUTO_architecture13 of FD_1801 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1546 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1546);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1800 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1800;

architecture SYN_PLUTO_architecture14 of FD_1800 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1547 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1547);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1799 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1799;

architecture SYN_PLUTO_architecture15 of FD_1799 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1548 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1548);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1798 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1798;

architecture SYN_PLUTO_architecture16 of FD_1798 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1549 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1549);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1797 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1797;

architecture SYN_PLUTO_architecture17 of FD_1797 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1550 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1550);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1796 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1796;

architecture SYN_PLUTO_architecture18 of FD_1796 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1551 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1551);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1795 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1795;

architecture SYN_PLUTO_architecture19 of FD_1795 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1552 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1552);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1794 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1794;

architecture SYN_PLUTO_architecture20 of FD_1794 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1553 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1553);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1793 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1793;

architecture SYN_PLUTO_architecture21 of FD_1793 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1554 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1554);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1792 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1792;

architecture SYN_PLUTO_architecture22 of FD_1792 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1555 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1555);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1791 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1791;

architecture SYN_PLUTO_architecture23 of FD_1791 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1556 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1556);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1790 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1790;

architecture SYN_PLUTO_architecture24 of FD_1790 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1557 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1557);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1789 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1789;

architecture SYN_PLUTO_architecture25 of FD_1789 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1558 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1558);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1788 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1788;

architecture SYN_PLUTO_architecture26 of FD_1788 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1559 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1559);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1787 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1787;

architecture SYN_PLUTO_architecture27 of FD_1787 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1560 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1560);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1786 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1786;

architecture SYN_PLUTO_architecture28 of FD_1786 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1561 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1561);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1785 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1785;

architecture SYN_PLUTO_architecture29 of FD_1785 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1562 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1562);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1784 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1784;

architecture SYN_PLUTO_architecture30 of FD_1784 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1563 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1563);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1783 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1783;

architecture SYN_PLUTO_architecture31 of FD_1783 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1564 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1564);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1782 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1782;

architecture SYN_PLUTO of FD_1782 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1565 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1565);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1781 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1781;

architecture SYN_PLUTO_architecture of FD_1781 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1566 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1566);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1780 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1780;

architecture SYN_PLUTO_architecture2 of FD_1780 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1567 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1567);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1779 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1779;

architecture SYN_PLUTO_architecture3 of FD_1779 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1568 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1568);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1778 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1778;

architecture SYN_PLUTO_architecture4 of FD_1778 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1569 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1569);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1777 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1777;

architecture SYN_PLUTO_architecture5 of FD_1777 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1570 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1570);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1776 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1776;

architecture SYN_PLUTO_architecture6 of FD_1776 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1571 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1571);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1775 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1775;

architecture SYN_PLUTO_architecture7 of FD_1775 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1572 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1572);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1774 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1774;

architecture SYN_PLUTO_architecture8 of FD_1774 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1573 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1573);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1773 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1773;

architecture SYN_PLUTO_architecture9 of FD_1773 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1574 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1574);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1772 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1772;

architecture SYN_PLUTO_architecture10 of FD_1772 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1575 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1575);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1771 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1771;

architecture SYN_PLUTO_architecture11 of FD_1771 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1576 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1576);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1770 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1770;

architecture SYN_PLUTO_architecture12 of FD_1770 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1577 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1577);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1769 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1769;

architecture SYN_PLUTO_architecture13 of FD_1769 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1578 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1578);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1768 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1768;

architecture SYN_PLUTO_architecture14 of FD_1768 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1579 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1579);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1767 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1767;

architecture SYN_PLUTO_architecture15 of FD_1767 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1580 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1580);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1766 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1766;

architecture SYN_PLUTO_architecture16 of FD_1766 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1581 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1581);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1765 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1765;

architecture SYN_PLUTO_architecture17 of FD_1765 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1582 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1582);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1764 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1764;

architecture SYN_PLUTO_architecture18 of FD_1764 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1583 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1583);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1763 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1763;

architecture SYN_PLUTO_architecture19 of FD_1763 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1584 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1584);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1762 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1762;

architecture SYN_PLUTO_architecture20 of FD_1762 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1585 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1585);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1761 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1761;

architecture SYN_PLUTO_architecture21 of FD_1761 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1586 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1586);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1760 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1760;

architecture SYN_PLUTO_architecture22 of FD_1760 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1587 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1587);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1759 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1759;

architecture SYN_PLUTO_architecture23 of FD_1759 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1588 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1588);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1758 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1758;

architecture SYN_PLUTO_architecture24 of FD_1758 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1589 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1589);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1757 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1757;

architecture SYN_PLUTO_architecture25 of FD_1757 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1590 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1590);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1756 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1756;

architecture SYN_PLUTO_architecture26 of FD_1756 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1591 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1591);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1755 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1755;

architecture SYN_PLUTO_architecture27 of FD_1755 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1592 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1592);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1754 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1754;

architecture SYN_PLUTO_architecture28 of FD_1754 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1593 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1593);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1753 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1753;

architecture SYN_PLUTO_architecture29 of FD_1753 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1594 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1594);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1752 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1752;

architecture SYN_PLUTO_architecture30 of FD_1752 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1595 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1595);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1751 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1751;

architecture SYN_PLUTO_architecture31 of FD_1751 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1596 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1596);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1750 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1750;

architecture SYN_PLUTO of FD_1750 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1597 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1597);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1749 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1749;

architecture SYN_PLUTO of FD_1749 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1598 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1598);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1748 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1748;

architecture SYN_PLUTO of FD_1748 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1599 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1599);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1747 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1747;

architecture SYN_PLUTO of FD_1747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1600 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1600);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1746 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1746;

architecture SYN_PLUTO of FD_1746 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1601 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1601);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1745 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1745;

architecture SYN_PLUTO of FD_1745 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1602 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1602);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1744 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1744;

architecture SYN_PLUTO of FD_1744 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1603 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1603);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1743 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1743;

architecture SYN_PLUTO of FD_1743 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1604 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1604);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1742 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1742;

architecture SYN_PLUTO of FD_1742 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1605 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1605);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1741 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1741;

architecture SYN_PLUTO of FD_1741 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1606 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1606);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1740 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1740;

architecture SYN_PLUTO of FD_1740 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1607 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1607);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1739 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1739;

architecture SYN_PLUTO of FD_1739 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1608 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1608);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1738 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1738;

architecture SYN_PLUTO of FD_1738 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1609 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1609);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1737 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1737;

architecture SYN_PLUTO of FD_1737 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1610 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1610);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1736 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1736;

architecture SYN_PLUTO of FD_1736 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1611 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1611);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1735 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1735;

architecture SYN_PLUTO of FD_1735 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1612 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1612);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1734 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1734;

architecture SYN_PLUTO of FD_1734 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1613 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1613);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1733 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1733;

architecture SYN_PLUTO of FD_1733 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1614 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1614);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1732 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1732;

architecture SYN_PLUTO of FD_1732 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1615 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1615);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1731 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1731;

architecture SYN_PLUTO of FD_1731 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1616 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1616);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1730 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1730;

architecture SYN_PLUTO of FD_1730 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1617 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1617);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1729 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1729;

architecture SYN_PLUTO of FD_1729 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1618 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1618);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1728 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1728;

architecture SYN_PLUTO of FD_1728 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1619 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1619);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1727 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1727;

architecture SYN_PLUTO of FD_1727 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1620 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1620);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1726 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1726;

architecture SYN_PLUTO of FD_1726 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1621 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1621);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1725 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1725;

architecture SYN_PLUTO of FD_1725 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1622 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1622);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1724 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1724;

architecture SYN_PLUTO of FD_1724 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1623 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1623);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1723 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1723;

architecture SYN_PLUTO of FD_1723 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1624 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1624);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1722 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1722;

architecture SYN_PLUTO of FD_1722 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1625 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1625);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1721 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1721;

architecture SYN_PLUTO of FD_1721 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1626 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1626);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1720 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1720;

architecture SYN_PLUTO of FD_1720 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1627 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1627);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1719 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1719;

architecture SYN_PLUTO of FD_1719 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1628 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1628);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1718 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1718;

architecture SYN_PLUTO of FD_1718 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1629 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1629);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1717 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1717;

architecture SYN_PLUTO of FD_1717 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1630 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1630);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1716 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1716;

architecture SYN_PLUTO of FD_1716 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1631 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1631);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1715 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1715;

architecture SYN_PLUTO of FD_1715 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1632 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1632);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1714 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1714;

architecture SYN_PLUTO of FD_1714 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1633 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1633);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1713 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1713;

architecture SYN_PLUTO of FD_1713 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1634 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1634);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1712 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1712;

architecture SYN_PLUTO of FD_1712 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1635 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1635);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1711 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1711;

architecture SYN_PLUTO of FD_1711 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1636 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1636);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1710 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1710;

architecture SYN_PLUTO of FD_1710 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1637 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1637);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1709 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1709;

architecture SYN_PLUTO of FD_1709 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1638 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1638);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1708 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1708;

architecture SYN_PLUTO of FD_1708 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1639 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1639);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1707 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1707;

architecture SYN_PLUTO of FD_1707 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1640 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1640);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1706 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1706;

architecture SYN_PLUTO of FD_1706 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1641 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1641);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1705 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1705;

architecture SYN_PLUTO of FD_1705 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1642 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1642);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1704 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1704;

architecture SYN_PLUTO of FD_1704 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1643 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1643);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1703 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1703;

architecture SYN_PLUTO of FD_1703 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1644 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1644);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1702 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1702;

architecture SYN_PLUTO of FD_1702 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1645 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1645);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1701 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1701;

architecture SYN_PLUTO of FD_1701 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1646 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1646);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1700 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1700;

architecture SYN_PLUTO of FD_1700 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1647 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1647);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1699 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1699;

architecture SYN_PLUTO of FD_1699 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1648 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1648);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1698 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1698;

architecture SYN_PLUTO of FD_1698 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1649 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1649);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1697 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1697;

architecture SYN_PLUTO of FD_1697 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1650 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1650);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1696 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1696;

architecture SYN_PLUTO of FD_1696 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1651 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1651);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1695 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1695;

architecture SYN_PLUTO of FD_1695 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1652 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1652);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1694 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1694;

architecture SYN_PLUTO of FD_1694 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1653 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1653);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1693 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1693;

architecture SYN_PLUTO of FD_1693 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1654 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1654);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1692 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1692;

architecture SYN_PLUTO of FD_1692 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1655 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1655);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1691 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1691;

architecture SYN_PLUTO of FD_1691 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1656 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1656);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1690 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1690;

architecture SYN_PLUTO of FD_1690 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1657 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1657);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1689 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1689;

architecture SYN_PLUTO of FD_1689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1658 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1658);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1688 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1688;

architecture SYN_PLUTO of FD_1688 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1659 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1659);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1687 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1687;

architecture SYN_PLUTO of FD_1687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1660 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1660);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1686 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1686;

architecture SYN_PLUTO of FD_1686 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1661 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1661);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1685 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1685;

architecture SYN_PLUTO of FD_1685 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1662 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1662);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1684 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1684;

architecture SYN_PLUTO of FD_1684 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1663 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1663);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1683 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1683;

architecture SYN_PLUTO of FD_1683 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1664 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1664);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1682 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1682;

architecture SYN_PLUTO of FD_1682 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1665 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1665);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1681 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1681;

architecture SYN_PLUTO of FD_1681 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1666 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1666);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1680 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1680;

architecture SYN_PLUTO of FD_1680 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1667 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1667);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1679 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1679;

architecture SYN_PLUTO of FD_1679 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1668 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1668);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1678 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1678;

architecture SYN_PLUTO of FD_1678 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1669 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1669);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1677 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1677;

architecture SYN_PLUTO of FD_1677 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1670 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1670);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1676 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1676;

architecture SYN_PLUTO of FD_1676 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1671 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1671);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1675 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1675;

architecture SYN_PLUTO of FD_1675 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1672 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1672);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1674 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1674;

architecture SYN_PLUTO of FD_1674 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1673 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1673);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1673 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1673;

architecture SYN_PLUTO of FD_1673 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1674 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1674);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1672 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1672;

architecture SYN_PLUTO of FD_1672 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1675 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1675);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1671 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1671;

architecture SYN_PLUTO of FD_1671 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1676 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1676);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1670 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1670;

architecture SYN_PLUTO of FD_1670 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1677 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1677);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1669 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1669;

architecture SYN_PLUTO of FD_1669 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1678 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1678);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1668 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1668;

architecture SYN_PLUTO of FD_1668 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1679 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1679);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1667 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1667;

architecture SYN_PLUTO of FD_1667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1680 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1680);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1666 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1666;

architecture SYN_PLUTO of FD_1666 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1681 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1681);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1665 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1665;

architecture SYN_PLUTO of FD_1665 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1682 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1682);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1664 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1664;

architecture SYN_PLUTO of FD_1664 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1683 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1683);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1663 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1663;

architecture SYN_PLUTO of FD_1663 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1684 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1684);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1662 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1662;

architecture SYN_PLUTO of FD_1662 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1685 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1685);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1661 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1661;

architecture SYN_PLUTO of FD_1661 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1686 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1686);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1660 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1660;

architecture SYN_PLUTO of FD_1660 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1687 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1687);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1659 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1659;

architecture SYN_PLUTO of FD_1659 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1688 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1688);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1658 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1658;

architecture SYN_PLUTO of FD_1658 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1689 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1689);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1657 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1657;

architecture SYN_PLUTO of FD_1657 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1690 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1690);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1656 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1656;

architecture SYN_PLUTO of FD_1656 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1691 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1691);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1655 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1655;

architecture SYN_PLUTO of FD_1655 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1692 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1692);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1654 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1654;

architecture SYN_PLUTO of FD_1654 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1693 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1693);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1653 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1653;

architecture SYN_PLUTO of FD_1653 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1694 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1694);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1652 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1652;

architecture SYN_PLUTO of FD_1652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1695 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1695);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1651 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1651;

architecture SYN_PLUTO of FD_1651 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1696 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1696);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1650 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1650;

architecture SYN_PLUTO of FD_1650 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1697 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1697);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1649 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1649;

architecture SYN_PLUTO of FD_1649 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1698 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1698);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1648 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1648;

architecture SYN_PLUTO of FD_1648 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1699 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1699);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1647 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1647;

architecture SYN_PLUTO of FD_1647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1700 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1700);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1646 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1646;

architecture SYN_PLUTO of FD_1646 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1701 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1701);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1645 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1645;

architecture SYN_PLUTO of FD_1645 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1702 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1702);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1644 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1644;

architecture SYN_PLUTO of FD_1644 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1703 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1703);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1643 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1643;

architecture SYN_PLUTO of FD_1643 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1704 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1704);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1642 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1642;

architecture SYN_PLUTO of FD_1642 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1705 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1705);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1641 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1641;

architecture SYN_PLUTO of FD_1641 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1706 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1706);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1640 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1640;

architecture SYN_PLUTO of FD_1640 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1707 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1707);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1639 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1639;

architecture SYN_PLUTO of FD_1639 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1708 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1708);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1638 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1638;

architecture SYN_PLUTO of FD_1638 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1709 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1709);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1637 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1637;

architecture SYN_PLUTO of FD_1637 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1710 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1710);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1636 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1636;

architecture SYN_PLUTO of FD_1636 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1711 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1711);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1635 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1635;

architecture SYN_PLUTO of FD_1635 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1712 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1712);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1634 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1634;

architecture SYN_PLUTO of FD_1634 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1713 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1713);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1633 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1633;

architecture SYN_PLUTO of FD_1633 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1714 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1714);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1632 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1632;

architecture SYN_PLUTO of FD_1632 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1715 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1715);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1631 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1631;

architecture SYN_PLUTO of FD_1631 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1716 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1716);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1630 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1630;

architecture SYN_PLUTO of FD_1630 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1717 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1717);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1629 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1629;

architecture SYN_PLUTO of FD_1629 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1718 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1718);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1628 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1628;

architecture SYN_PLUTO of FD_1628 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1719 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1719);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1627 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1627;

architecture SYN_PLUTO of FD_1627 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1720 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1720);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1626 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1626;

architecture SYN_PLUTO of FD_1626 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1721 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1721);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1625 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1625;

architecture SYN_PLUTO of FD_1625 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1722 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1722);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1624 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1624;

architecture SYN_PLUTO of FD_1624 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1723 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1723);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1623 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1623;

architecture SYN_PLUTO of FD_1623 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1724 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1724);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1622 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1622;

architecture SYN_PLUTO of FD_1622 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1725 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1725);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1621 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1621;

architecture SYN_PLUTO of FD_1621 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1726 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1726);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1620 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1620;

architecture SYN_PLUTO of FD_1620 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1727 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1727);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1619 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1619;

architecture SYN_PLUTO of FD_1619 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1728 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1728);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1618 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1618;

architecture SYN_PLUTO of FD_1618 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1729 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1729);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1617 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1617;

architecture SYN_PLUTO of FD_1617 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1730 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1730);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1616 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1616;

architecture SYN_PLUTO of FD_1616 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1731 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1731);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1615 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1615;

architecture SYN_PLUTO of FD_1615 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1732 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1732);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1614 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1614;

architecture SYN_PLUTO of FD_1614 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1733 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1733);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1613 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1613;

architecture SYN_PLUTO of FD_1613 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1734 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1734);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1612 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1612;

architecture SYN_PLUTO of FD_1612 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1735 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1735);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1611 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1611;

architecture SYN_PLUTO of FD_1611 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1736 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1736);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1610 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1610;

architecture SYN_PLUTO of FD_1610 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1737 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1737);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1609 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1609;

architecture SYN_PLUTO of FD_1609 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1738 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1738);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1608 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1608;

architecture SYN_PLUTO of FD_1608 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1739 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1739);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1607 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1607;

architecture SYN_PLUTO of FD_1607 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1740 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1740);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1606 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1606;

architecture SYN_PLUTO of FD_1606 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1741 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1741);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1605 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1605;

architecture SYN_PLUTO of FD_1605 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1742 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1742);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1604 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1604;

architecture SYN_PLUTO of FD_1604 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1743 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1743);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1603 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1603;

architecture SYN_PLUTO of FD_1603 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1744 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1744);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1602 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1602;

architecture SYN_PLUTO of FD_1602 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1745 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1745);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1601 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1601;

architecture SYN_PLUTO of FD_1601 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1746 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1746);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1600 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1600;

architecture SYN_PLUTO of FD_1600 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1747 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1747);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1599 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1599;

architecture SYN_PLUTO of FD_1599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1748 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1748);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1598 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1598;

architecture SYN_PLUTO of FD_1598 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1749 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1749);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1597 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1597;

architecture SYN_PLUTO of FD_1597 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1750 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1750);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1596 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1596;

architecture SYN_PLUTO of FD_1596 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1751 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1751);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1595 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1595;

architecture SYN_PLUTO of FD_1595 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1752 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1752);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1594 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1594;

architecture SYN_PLUTO of FD_1594 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1753 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1753);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1593 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1593;

architecture SYN_PLUTO of FD_1593 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1754 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1754);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1592 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1592;

architecture SYN_PLUTO of FD_1592 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1755 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1755);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1591 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1591;

architecture SYN_PLUTO of FD_1591 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1756 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1756);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1590 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1590;

architecture SYN_PLUTO of FD_1590 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1757 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1757);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1589 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1589;

architecture SYN_PLUTO of FD_1589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1758 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1758);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1588 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1588;

architecture SYN_PLUTO of FD_1588 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1759 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1759);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1587 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1587;

architecture SYN_PLUTO of FD_1587 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1760 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1760);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1586 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1586;

architecture SYN_PLUTO of FD_1586 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1761 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1761);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1585 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1585;

architecture SYN_PLUTO of FD_1585 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1762 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1762);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1584 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1584;

architecture SYN_PLUTO of FD_1584 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1763 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1763);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1583 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1583;

architecture SYN_PLUTO of FD_1583 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1764 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1764);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1582 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1582;

architecture SYN_PLUTO of FD_1582 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1765 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1765);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1581 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1581;

architecture SYN_PLUTO of FD_1581 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1766 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1766);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1580 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1580;

architecture SYN_PLUTO of FD_1580 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1767 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1767);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1579 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1579;

architecture SYN_PLUTO of FD_1579 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1768 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1768);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1578 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1578;

architecture SYN_PLUTO of FD_1578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1769 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1769);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1577 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1577;

architecture SYN_PLUTO of FD_1577 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1770 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1770);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1576 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1576;

architecture SYN_PLUTO of FD_1576 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1771 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1771);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1575 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1575;

architecture SYN_PLUTO of FD_1575 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1772 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1772);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1574 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1574;

architecture SYN_PLUTO of FD_1574 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1773 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1773);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1573 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1573;

architecture SYN_PLUTO of FD_1573 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1774 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1774);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1572 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1572;

architecture SYN_PLUTO of FD_1572 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1775 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1775);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1571 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1571;

architecture SYN_PLUTO of FD_1571 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1776 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1776);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1570 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1570;

architecture SYN_PLUTO of FD_1570 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1777 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1777);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1569 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1569;

architecture SYN_PLUTO of FD_1569 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1778 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1778);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1568 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1568;

architecture SYN_PLUTO of FD_1568 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1779 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1779);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1567 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1567;

architecture SYN_PLUTO of FD_1567 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1780 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1780);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1566 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1566;

architecture SYN_PLUTO of FD_1566 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1781 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1781);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1565 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1565;

architecture SYN_PLUTO of FD_1565 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1782 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1782);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1564 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1564;

architecture SYN_PLUTO of FD_1564 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1783 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1783);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1563 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1563;

architecture SYN_PLUTO of FD_1563 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1784 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1784);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1562 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1562;

architecture SYN_PLUTO of FD_1562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1785 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1785);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1561 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1561;

architecture SYN_PLUTO of FD_1561 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1786 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1786);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1560 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1560;

architecture SYN_PLUTO of FD_1560 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1787 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1787);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1559 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1559;

architecture SYN_PLUTO of FD_1559 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1788 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1788);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1558 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1558;

architecture SYN_PLUTO of FD_1558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1789 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1789);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1557 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1557;

architecture SYN_PLUTO of FD_1557 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1790 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1790);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1556 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1556;

architecture SYN_PLUTO of FD_1556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1791 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1791);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1555 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1555;

architecture SYN_PLUTO of FD_1555 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1792 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1792);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1554 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1554;

architecture SYN_PLUTO of FD_1554 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1793 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1793);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1553 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1553;

architecture SYN_PLUTO of FD_1553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1794 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1794);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1552 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1552;

architecture SYN_PLUTO of FD_1552 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1795 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1795);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1551 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1551;

architecture SYN_PLUTO of FD_1551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1796 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1796);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1550 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1550;

architecture SYN_PLUTO of FD_1550 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1797 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1797);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1549 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1549;

architecture SYN_PLUTO of FD_1549 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1798 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1798);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1548 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1548;

architecture SYN_PLUTO of FD_1548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1799 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1799);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1547 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1547;

architecture SYN_PLUTO of FD_1547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1800 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1800);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1546 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1546;

architecture SYN_PLUTO of FD_1546 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1801 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1801);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1545 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1545;

architecture SYN_PLUTO of FD_1545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1802 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1802);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1544 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1544;

architecture SYN_PLUTO of FD_1544 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1803 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1803);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1543 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1543;

architecture SYN_PLUTO of FD_1543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1804 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1804);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1542 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1542;

architecture SYN_PLUTO of FD_1542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1805 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1805);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1541 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1541;

architecture SYN_PLUTO of FD_1541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1806 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1806);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1540 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1540;

architecture SYN_PLUTO of FD_1540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1807 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1807);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1539 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1539;

architecture SYN_PLUTO of FD_1539 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1808 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1808);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1538 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1538;

architecture SYN_PLUTO of FD_1538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1809 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1809);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1537 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1537;

architecture SYN_PLUTO of FD_1537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1810 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1810);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1536 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1536;

architecture SYN_PLUTO of FD_1536 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1811 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1811);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1535 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1535;

architecture SYN_PLUTO of FD_1535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1812 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1812);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1534 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1534;

architecture SYN_PLUTO of FD_1534 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1813 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1813);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1533 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1533;

architecture SYN_PLUTO of FD_1533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1814 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1814);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1532 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1532;

architecture SYN_PLUTO of FD_1532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1815 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1815);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1531 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1531;

architecture SYN_PLUTO of FD_1531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1816 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1816);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1530 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1530;

architecture SYN_PLUTO of FD_1530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1817 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1817);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1529 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1529;

architecture SYN_PLUTO of FD_1529 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1818 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1818);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1528 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1528;

architecture SYN_PLUTO of FD_1528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1819 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1819);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1527 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1527;

architecture SYN_PLUTO of FD_1527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1820 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1820);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1526 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1526;

architecture SYN_PLUTO of FD_1526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1821 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1821);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1525 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1525;

architecture SYN_PLUTO of FD_1525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1822 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1822);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1524 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1524;

architecture SYN_PLUTO of FD_1524 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1823 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1823);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1523 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1523;

architecture SYN_PLUTO of FD_1523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1824 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1824);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1522 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1522;

architecture SYN_PLUTO of FD_1522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1825 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1825);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1521 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1521;

architecture SYN_PLUTO of FD_1521 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1826 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1826);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1520 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1520;

architecture SYN_PLUTO of FD_1520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1827 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1827);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1519 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1519;

architecture SYN_PLUTO of FD_1519 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1828 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1828);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1518 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1518;

architecture SYN_PLUTO of FD_1518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1829 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1829);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1517 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1517;

architecture SYN_PLUTO of FD_1517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1830 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1830);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1516 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1516;

architecture SYN_PLUTO of FD_1516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1831 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1831);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1515 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1515;

architecture SYN_PLUTO of FD_1515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1832 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1832);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1514 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1514;

architecture SYN_PLUTO of FD_1514 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1833 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1833);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1513 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1513;

architecture SYN_PLUTO of FD_1513 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1834 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1834);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1512 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1512;

architecture SYN_PLUTO of FD_1512 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1835 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1835);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1511 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1511;

architecture SYN_PLUTO of FD_1511 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1836 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1836);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1510 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1510;

architecture SYN_PLUTO of FD_1510 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1837 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1837);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1509 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1509;

architecture SYN_PLUTO of FD_1509 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1838 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1838);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1508 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1508;

architecture SYN_PLUTO of FD_1508 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1839 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1839);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1507 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1507;

architecture SYN_PLUTO of FD_1507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1840 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1840);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1506 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1506;

architecture SYN_PLUTO of FD_1506 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1841 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1841);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1505 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1505;

architecture SYN_PLUTO of FD_1505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1842 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1842);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1504 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1504;

architecture SYN_PLUTO of FD_1504 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1843 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1843);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1503 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1503;

architecture SYN_PLUTO of FD_1503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1844 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1844);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1502 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1502;

architecture SYN_PLUTO of FD_1502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1845 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1845);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1501 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1501;

architecture SYN_PLUTO of FD_1501 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1846 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1846);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1500 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1500;

architecture SYN_PLUTO_architecture of FD_1500 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1847 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1847);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1499 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1499;

architecture SYN_PLUTO_architecture2 of FD_1499 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1848 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1848);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1498 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1498;

architecture SYN_PLUTO_architecture3 of FD_1498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1849 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1849);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1497 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1497;

architecture SYN_PLUTO_architecture4 of FD_1497 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1850 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1850);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1496 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1496;

architecture SYN_PLUTO_architecture5 of FD_1496 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1851 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1851);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1495 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1495;

architecture SYN_PLUTO_architecture6 of FD_1495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1852 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1852);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1494 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1494;

architecture SYN_PLUTO_architecture7 of FD_1494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1853 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1853);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1493 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1493;

architecture SYN_PLUTO_architecture8 of FD_1493 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1854 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1854);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1492 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1492;

architecture SYN_PLUTO_architecture9 of FD_1492 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1855 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1855);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1491 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1491;

architecture SYN_PLUTO_architecture10 of FD_1491 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1856 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1856);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1490 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1490;

architecture SYN_PLUTO_architecture11 of FD_1490 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1857 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1857);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1489 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1489;

architecture SYN_PLUTO_architecture12 of FD_1489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1858 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1858);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1488 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1488;

architecture SYN_PLUTO_architecture13 of FD_1488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1859 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1859);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1487 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1487;

architecture SYN_PLUTO_architecture14 of FD_1487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1860 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1860);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1486 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1486;

architecture SYN_PLUTO_architecture15 of FD_1486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1861 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1861);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1485 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1485;

architecture SYN_PLUTO_architecture16 of FD_1485 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1862 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1862);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1484 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1484;

architecture SYN_PLUTO_architecture17 of FD_1484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1863 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1863);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1483 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1483;

architecture SYN_PLUTO_architecture18 of FD_1483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1864 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1864);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1482 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1482;

architecture SYN_PLUTO_architecture19 of FD_1482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1865 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1865);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1481 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1481;

architecture SYN_PLUTO_architecture20 of FD_1481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1866 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1866);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1480 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1480;

architecture SYN_PLUTO_architecture21 of FD_1480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1867 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1867);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1479 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1479;

architecture SYN_PLUTO_architecture22 of FD_1479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1868 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1868);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1478 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1478;

architecture SYN_PLUTO_architecture23 of FD_1478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1869 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1869);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1477 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1477;

architecture SYN_PLUTO_architecture24 of FD_1477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1870 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1870);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1476 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1476;

architecture SYN_PLUTO_architecture25 of FD_1476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1871 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1871);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1475 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1475;

architecture SYN_PLUTO_architecture26 of FD_1475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1872 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1872);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1474 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1474;

architecture SYN_PLUTO_architecture27 of FD_1474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1873 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1873);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1473 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1473;

architecture SYN_PLUTO_architecture28 of FD_1473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1874 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1874);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1472 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1472;

architecture SYN_PLUTO_architecture29 of FD_1472 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1875 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1875);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1471 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1471;

architecture SYN_PLUTO_architecture30 of FD_1471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1876 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1876);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1470 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1470;

architecture SYN_PLUTO_architecture31 of FD_1470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1877 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1877);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1469 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1469;

architecture SYN_PLUTO of FD_1469 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1878 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1878);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1468 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1468;

architecture SYN_PLUTO_architecture of FD_1468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1879 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1879);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1467 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1467;

architecture SYN_PLUTO_architecture2 of FD_1467 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1880 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1880);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1466 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1466;

architecture SYN_PLUTO_architecture3 of FD_1466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1881 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1881);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1465 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1465;

architecture SYN_PLUTO_architecture4 of FD_1465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1882 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1882);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1464 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1464;

architecture SYN_PLUTO_architecture5 of FD_1464 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1883 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1883);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1463 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1463;

architecture SYN_PLUTO_architecture6 of FD_1463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1884 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1884);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1462 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1462;

architecture SYN_PLUTO_architecture7 of FD_1462 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1885 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1885);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1461 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1461;

architecture SYN_PLUTO_architecture8 of FD_1461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1886 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1886);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1460 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1460;

architecture SYN_PLUTO_architecture9 of FD_1460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1887 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1887);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1459 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1459;

architecture SYN_PLUTO_architecture10 of FD_1459 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1888 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1888);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1458 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1458;

architecture SYN_PLUTO_architecture11 of FD_1458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1889 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1889);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1457 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1457;

architecture SYN_PLUTO_architecture12 of FD_1457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1890 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1890);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1456 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1456;

architecture SYN_PLUTO_architecture13 of FD_1456 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1891 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1891);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1455 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1455;

architecture SYN_PLUTO_architecture14 of FD_1455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1892 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1892);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1454 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1454;

architecture SYN_PLUTO_architecture15 of FD_1454 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1893 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1893);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1453 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1453;

architecture SYN_PLUTO_architecture16 of FD_1453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1894 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1894);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1452 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1452;

architecture SYN_PLUTO_architecture17 of FD_1452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1895 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1895);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1451 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1451;

architecture SYN_PLUTO_architecture18 of FD_1451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1896 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1896);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1450 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1450;

architecture SYN_PLUTO_architecture19 of FD_1450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1897 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1897);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1449 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1449;

architecture SYN_PLUTO_architecture20 of FD_1449 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1898 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1898);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1448 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1448;

architecture SYN_PLUTO_architecture21 of FD_1448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1899 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1899);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1447 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1447;

architecture SYN_PLUTO_architecture22 of FD_1447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1900 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1900);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1446 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1446;

architecture SYN_PLUTO_architecture23 of FD_1446 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1901 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1901);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1445 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1445;

architecture SYN_PLUTO_architecture24 of FD_1445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1902 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1902);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1444 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1444;

architecture SYN_PLUTO_architecture25 of FD_1444 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1903 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1903);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1443 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1443;

architecture SYN_PLUTO_architecture26 of FD_1443 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1904 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1904);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1442 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1442;

architecture SYN_PLUTO_architecture27 of FD_1442 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1905 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1905);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1441 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1441;

architecture SYN_PLUTO_architecture28 of FD_1441 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1906 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1906);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1440 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1440;

architecture SYN_PLUTO_architecture29 of FD_1440 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1907 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1907);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1439 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1439;

architecture SYN_PLUTO_architecture30 of FD_1439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1908 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1908);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1438 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1438;

architecture SYN_PLUTO_architecture31 of FD_1438 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1909 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1909);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1437 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1437;

architecture SYN_PLUTO_architecture32 of FD_1437 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1910 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1910);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1436 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1436;

architecture SYN_PLUTO_architecture33 of FD_1436 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1911 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1911);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1435 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1435;

architecture SYN_PLUTO_architecture34 of FD_1435 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1912 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1912);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1434 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1434;

architecture SYN_PLUTO_architecture35 of FD_1434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1913 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1913);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1433 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1433;

architecture SYN_PLUTO_architecture36 of FD_1433 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1914 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1914);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1432 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1432;

architecture SYN_PLUTO_architecture37 of FD_1432 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1915 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1915);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1431 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1431;

architecture SYN_PLUTO_architecture38 of FD_1431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1916 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1916);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1430 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1430;

architecture SYN_PLUTO_architecture39 of FD_1430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1917 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1917);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1429 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1429;

architecture SYN_PLUTO_architecture40 of FD_1429 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1918 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1918);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1428 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1428;

architecture SYN_PLUTO_architecture41 of FD_1428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1919 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1919);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1427 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1427;

architecture SYN_PLUTO_architecture42 of FD_1427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1920 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1920);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1426 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1426;

architecture SYN_PLUTO_architecture43 of FD_1426 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1921 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1921);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1425 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1425;

architecture SYN_PLUTO_architecture44 of FD_1425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1922 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1922);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1424 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1424;

architecture SYN_PLUTO_architecture45 of FD_1424 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1923 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1923);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1423 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1423;

architecture SYN_PLUTO_architecture46 of FD_1423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1924 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1924);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1422 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1422;

architecture SYN_PLUTO_architecture47 of FD_1422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1925 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1925);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1421 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1421;

architecture SYN_PLUTO_architecture48 of FD_1421 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1926 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1926);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1420 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1420;

architecture SYN_PLUTO_architecture49 of FD_1420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1927 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1927);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1419 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1419;

architecture SYN_PLUTO_architecture50 of FD_1419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1928 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1928);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1418 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1418;

architecture SYN_PLUTO_architecture51 of FD_1418 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1929 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1929);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1417 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1417;

architecture SYN_PLUTO_architecture52 of FD_1417 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1930 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1930);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1416 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1416;

architecture SYN_PLUTO_architecture53 of FD_1416 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1931 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1931);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1415 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1415;

architecture SYN_PLUTO_architecture54 of FD_1415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1932 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1932);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1414 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1414;

architecture SYN_PLUTO_architecture55 of FD_1414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1933 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1933);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1413 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1413;

architecture SYN_PLUTO_architecture56 of FD_1413 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1934 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1934);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1412 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1412;

architecture SYN_PLUTO_architecture57 of FD_1412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1935 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1935);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1411 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1411;

architecture SYN_PLUTO_architecture58 of FD_1411 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1936 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1936);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1410 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1410;

architecture SYN_PLUTO_architecture59 of FD_1410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1937 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1937);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1409 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1409;

architecture SYN_PLUTO_architecture60 of FD_1409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1938 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1938);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1408 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1408;

architecture SYN_PLUTO_architecture61 of FD_1408 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1939 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1939);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1407 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1407;

architecture SYN_PLUTO_architecture62 of FD_1407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1940 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1940);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1406 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1406;

architecture SYN_PLUTO_architecture63 of FD_1406 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1941 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1941);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1405 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1405;

architecture SYN_PLUTO_architecture64 of FD_1405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1942 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1942);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1404 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1404;

architecture SYN_PLUTO_architecture65 of FD_1404 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1943 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1943);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1403 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1403;

architecture SYN_PLUTO_architecture66 of FD_1403 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1944 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1944);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1402 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1402;

architecture SYN_PLUTO_architecture67 of FD_1402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1945 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1945);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1401 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1401;

architecture SYN_PLUTO_architecture68 of FD_1401 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1946 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1946);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1400 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1400;

architecture SYN_PLUTO_architecture69 of FD_1400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1947 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1947);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1399 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1399;

architecture SYN_PLUTO_architecture70 of FD_1399 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1948 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1948);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1398 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1398;

architecture SYN_PLUTO_architecture71 of FD_1398 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1949 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1949);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1397 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1397;

architecture SYN_PLUTO_architecture72 of FD_1397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1950 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1950);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1396 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1396;

architecture SYN_PLUTO_architecture73 of FD_1396 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1951 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1951);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1395 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1395;

architecture SYN_PLUTO_architecture74 of FD_1395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1952 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1952);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1394 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1394;

architecture SYN_PLUTO_architecture75 of FD_1394 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1953 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1953);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1393 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1393;

architecture SYN_PLUTO_architecture76 of FD_1393 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1954 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1954);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1392 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1392;

architecture SYN_PLUTO_architecture77 of FD_1392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1955 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1955);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1391 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1391;

architecture SYN_PLUTO_architecture78 of FD_1391 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1956 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1956);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1390 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1390;

architecture SYN_PLUTO_architecture79 of FD_1390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1957 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1957);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1389 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1389;

architecture SYN_PLUTO_architecture80 of FD_1389 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1958 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1958);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1388 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1388;

architecture SYN_PLUTO_architecture81 of FD_1388 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1959 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1959);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1387 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1387;

architecture SYN_PLUTO_architecture82 of FD_1387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1960 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1960);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1386 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1386;

architecture SYN_PLUTO_architecture83 of FD_1386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1961 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1961);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1385 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1385;

architecture SYN_PLUTO_architecture84 of FD_1385 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1962 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1962);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1384 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1384;

architecture SYN_PLUTO_architecture85 of FD_1384 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1963 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1963);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1383 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1383;

architecture SYN_PLUTO_architecture86 of FD_1383 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1964 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1964);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1382 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1382;

architecture SYN_PLUTO_architecture87 of FD_1382 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1965 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1965);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1381 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1381;

architecture SYN_PLUTO_architecture88 of FD_1381 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1966 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1966);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1380 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1380;

architecture SYN_PLUTO_architecture89 of FD_1380 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1967 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1967);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1379 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1379;

architecture SYN_PLUTO_architecture90 of FD_1379 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1968 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1968);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1378 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1378;

architecture SYN_PLUTO_architecture91 of FD_1378 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1969 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1969);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1377 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1377;

architecture SYN_PLUTO_architecture92 of FD_1377 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1970 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1970);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1376 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1376;

architecture SYN_PLUTO_architecture93 of FD_1376 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1971 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1971);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1375 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1375;

architecture SYN_PLUTO_architecture94 of FD_1375 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1972 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1972);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1374 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1374;

architecture SYN_PLUTO_architecture95 of FD_1374 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1973 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1973);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1373 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1373;

architecture SYN_PLUTO_architecture96 of FD_1373 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1974 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1974);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1372 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1372;

architecture SYN_PLUTO_architecture97 of FD_1372 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1975 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1975);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1371 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1371;

architecture SYN_PLUTO_architecture98 of FD_1371 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1976 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1976);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1370 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1370;

architecture SYN_PLUTO_architecture99 of FD_1370 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1977 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1977);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1369 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1369;

architecture SYN_PLUTO_architecture100 of FD_1369 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1978 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1978);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1368 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1368;

architecture SYN_PLUTO_architecture101 of FD_1368 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1979 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1979);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1367 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1367;

architecture SYN_PLUTO_architecture102 of FD_1367 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1980 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1980);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1366 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1366;

architecture SYN_PLUTO_architecture103 of FD_1366 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1981 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1981);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1365 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1365;

architecture SYN_PLUTO_architecture104 of FD_1365 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1982 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1982);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1364 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1364;

architecture SYN_PLUTO_architecture105 of FD_1364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1983 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1983);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1363 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1363;

architecture SYN_PLUTO_architecture106 of FD_1363 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1984 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1984);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1362 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1362;

architecture SYN_PLUTO_architecture107 of FD_1362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1985 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1985);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1361 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1361;

architecture SYN_PLUTO_architecture108 of FD_1361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1986 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1986);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1360 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1360;

architecture SYN_PLUTO_architecture109 of FD_1360 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1987 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1987);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1359 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1359;

architecture SYN_PLUTO_architecture110 of FD_1359 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1988 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1988);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1358 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1358;

architecture SYN_PLUTO_architecture111 of FD_1358 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1989 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1989);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1357 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1357;

architecture SYN_PLUTO_architecture112 of FD_1357 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1990 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1990);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1356 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1356;

architecture SYN_PLUTO_architecture113 of FD_1356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1991 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1991);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1355 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1355;

architecture SYN_PLUTO_architecture114 of FD_1355 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1992 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1992);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1354 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1354;

architecture SYN_PLUTO_architecture115 of FD_1354 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1993 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1993);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1353 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1353;

architecture SYN_PLUTO_architecture116 of FD_1353 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1994 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1994);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1352 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1352;

architecture SYN_PLUTO_architecture117 of FD_1352 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1995 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1995);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1351 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1351;

architecture SYN_PLUTO_architecture118 of FD_1351 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1996 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1996);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1350 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1350;

architecture SYN_PLUTO_architecture119 of FD_1350 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1997 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1997);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1349 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1349;

architecture SYN_PLUTO_architecture120 of FD_1349 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1998 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1998);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1348 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1348;

architecture SYN_PLUTO_architecture121 of FD_1348 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_1999 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_1999);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1347 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1347;

architecture SYN_PLUTO_architecture122 of FD_1347 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2000 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2000);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1346 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1346;

architecture SYN_PLUTO_architecture123 of FD_1346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2001 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2001);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1345 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1345;

architecture SYN_PLUTO_architecture124 of FD_1345 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2002 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2002);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1344 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1344;

architecture SYN_PLUTO_architecture125 of FD_1344 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2003 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2003);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1343 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1343;

architecture SYN_PLUTO_architecture126 of FD_1343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2004 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2004);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1342 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1342;

architecture SYN_PLUTO_architecture127 of FD_1342 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2005 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2005);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1341 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1341;

architecture SYN_PLUTO_architecture128 of FD_1341 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2006 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2006);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1340 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1340;

architecture SYN_PLUTO_architecture129 of FD_1340 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2007 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2007);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1339 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1339;

architecture SYN_PLUTO_architecture130 of FD_1339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2008 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2008);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1338 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1338;

architecture SYN_PLUTO_architecture131 of FD_1338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2009 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2009);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1337 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1337;

architecture SYN_PLUTO_architecture132 of FD_1337 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2010 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2010);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1336 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1336;

architecture SYN_PLUTO_architecture133 of FD_1336 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2011 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2011);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1335 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1335;

architecture SYN_PLUTO_architecture134 of FD_1335 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2012 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2012);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1334 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1334;

architecture SYN_PLUTO_architecture135 of FD_1334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2013 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2013);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1333 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1333;

architecture SYN_PLUTO_architecture136 of FD_1333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2014 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2014);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1332 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1332;

architecture SYN_PLUTO_architecture137 of FD_1332 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2015 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2015);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1331 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1331;

architecture SYN_PLUTO_architecture138 of FD_1331 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2016 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2016);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1330 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1330;

architecture SYN_PLUTO_architecture139 of FD_1330 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2017 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2017);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1329 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1329;

architecture SYN_PLUTO_architecture140 of FD_1329 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2018 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2018);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1328 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1328;

architecture SYN_PLUTO_architecture141 of FD_1328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2019 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2019);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1327 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1327;

architecture SYN_PLUTO_architecture142 of FD_1327 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2020 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2020);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1326 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1326;

architecture SYN_PLUTO_architecture143 of FD_1326 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2021 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2021);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture143;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1325 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1325;

architecture SYN_PLUTO_architecture144 of FD_1325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2022 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2022);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture144;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1324 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1324;

architecture SYN_PLUTO_architecture145 of FD_1324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2023 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2023);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture145;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1323 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1323;

architecture SYN_PLUTO_architecture146 of FD_1323 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2024 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2024);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture146;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1322 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1322;

architecture SYN_PLUTO_architecture147 of FD_1322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2025 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2025);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture147;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1321 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1321;

architecture SYN_PLUTO_architecture148 of FD_1321 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2026 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2026);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture148;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1320 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1320;

architecture SYN_PLUTO_architecture149 of FD_1320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2027 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2027);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture149;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1319 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1319;

architecture SYN_PLUTO_architecture150 of FD_1319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2028 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2028);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture150;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1318 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1318;

architecture SYN_PLUTO_architecture151 of FD_1318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2029 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2029);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture151;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1317 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1317;

architecture SYN_PLUTO_architecture152 of FD_1317 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2030 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2030);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture152;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1316 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1316;

architecture SYN_PLUTO_architecture153 of FD_1316 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2031 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2031);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture153;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1315 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1315;

architecture SYN_PLUTO_architecture154 of FD_1315 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2032 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2032);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture154;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1314 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1314;

architecture SYN_PLUTO_architecture155 of FD_1314 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2033 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2033);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture155;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1313 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1313;

architecture SYN_PLUTO_architecture156 of FD_1313 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2034 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2034);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture156;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1312 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1312;

architecture SYN_PLUTO_architecture157 of FD_1312 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2035 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2035);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture157;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1311 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1311;

architecture SYN_PLUTO_architecture158 of FD_1311 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2036 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2036);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture158;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1310 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1310;

architecture SYN_PLUTO_architecture159 of FD_1310 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2037 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2037);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture159;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1309 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1309;

architecture SYN_PLUTO_architecture160 of FD_1309 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2038 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2038);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture160;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1308 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1308;

architecture SYN_PLUTO_architecture161 of FD_1308 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2039 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2039);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture161;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1307 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1307;

architecture SYN_PLUTO_architecture162 of FD_1307 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2040 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2040);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture162;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1306 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1306;

architecture SYN_PLUTO_architecture163 of FD_1306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2041 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2041);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture163;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1305 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1305;

architecture SYN_PLUTO_architecture164 of FD_1305 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2042 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2042);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture164;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1304 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1304;

architecture SYN_PLUTO_architecture165 of FD_1304 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2043 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2043);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture165;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1303 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1303;

architecture SYN_PLUTO_architecture166 of FD_1303 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2044 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2044);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture166;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1302 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1302;

architecture SYN_PLUTO_architecture167 of FD_1302 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2045 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2045);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture167;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1301 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1301;

architecture SYN_PLUTO_architecture168 of FD_1301 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2046 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2046);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture168;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1300 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1300;

architecture SYN_PLUTO_architecture169 of FD_1300 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2047 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2047);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture169;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1299 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1299;

architecture SYN_PLUTO_architecture170 of FD_1299 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2048 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2048);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture170;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1298 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1298;

architecture SYN_PLUTO_architecture171 of FD_1298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2049 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2049);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture171;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1297 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1297;

architecture SYN_PLUTO_architecture172 of FD_1297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2050 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2050);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture172;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1296 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1296;

architecture SYN_PLUTO_architecture173 of FD_1296 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2051 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2051);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture173;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1295 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1295;

architecture SYN_PLUTO_architecture174 of FD_1295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2052 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2052);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture174;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1294 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1294;

architecture SYN_PLUTO_architecture175 of FD_1294 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2053 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2053);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture175;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1293 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1293;

architecture SYN_PLUTO_architecture176 of FD_1293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2054 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2054);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture176;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1292 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1292;

architecture SYN_PLUTO_architecture177 of FD_1292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2055 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2055);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture177;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1291 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1291;

architecture SYN_PLUTO_architecture178 of FD_1291 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2056 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2056);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture178;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1290 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1290;

architecture SYN_PLUTO_architecture179 of FD_1290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2057 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2057);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture179;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1289 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1289;

architecture SYN_PLUTO_architecture180 of FD_1289 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2058 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2058);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture180;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1288 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1288;

architecture SYN_PLUTO_architecture181 of FD_1288 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2059 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2059);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture181;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1287 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1287;

architecture SYN_PLUTO_architecture182 of FD_1287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2060 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2060);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture182;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1286 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1286;

architecture SYN_PLUTO_architecture183 of FD_1286 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2061 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2061);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture183;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1285 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1285;

architecture SYN_PLUTO_architecture184 of FD_1285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2062 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2062);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture184;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1284 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1284;

architecture SYN_PLUTO_architecture185 of FD_1284 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2063 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2063);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture185;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1283 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1283;

architecture SYN_PLUTO_architecture186 of FD_1283 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2064 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2064);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture186;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1282 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1282;

architecture SYN_PLUTO_architecture187 of FD_1282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2065 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2065);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture187;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1281 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1281;

architecture SYN_PLUTO_architecture188 of FD_1281 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2066 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2066);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture188;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1280 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1280;

architecture SYN_PLUTO_architecture189 of FD_1280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2067 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2067);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture189;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1279 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1279;

architecture SYN_PLUTO_architecture190 of FD_1279 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2068 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2068);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture190;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1278 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1278;

architecture SYN_PLUTO_architecture191 of FD_1278 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2069 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2069);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture191;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1277 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1277;

architecture SYN_PLUTO_architecture192 of FD_1277 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2070 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2070);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture192;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1276 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1276;

architecture SYN_PLUTO_architecture193 of FD_1276 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2071 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2071);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture193;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1275 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1275;

architecture SYN_PLUTO_architecture194 of FD_1275 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2072 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2072);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture194;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1274 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1274;

architecture SYN_PLUTO_architecture195 of FD_1274 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2073 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2073);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture195;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1273 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1273;

architecture SYN_PLUTO_architecture196 of FD_1273 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2074 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2074);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture196;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1272 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1272;

architecture SYN_PLUTO_architecture197 of FD_1272 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2075 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2075);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture197;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1271 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1271;

architecture SYN_PLUTO_architecture198 of FD_1271 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2076 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2076);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture198;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1270 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1270;

architecture SYN_PLUTO_architecture199 of FD_1270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2077 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2077);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture199;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1269 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1269;

architecture SYN_PLUTO_architecture200 of FD_1269 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2078 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2078);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture200;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1268 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1268;

architecture SYN_PLUTO_architecture201 of FD_1268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2079 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2079);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture201;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1267 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1267;

architecture SYN_PLUTO_architecture202 of FD_1267 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2080 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2080);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture202;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1266 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1266;

architecture SYN_PLUTO_architecture203 of FD_1266 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2081 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2081);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture203;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1265 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1265;

architecture SYN_PLUTO_architecture204 of FD_1265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2082 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2082);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture204;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1264 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1264;

architecture SYN_PLUTO_architecture205 of FD_1264 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2083 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2083);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture205;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1263 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1263;

architecture SYN_PLUTO_architecture206 of FD_1263 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2084 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2084);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture206;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1262 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1262;

architecture SYN_PLUTO_architecture207 of FD_1262 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2085 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2085);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture207;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1261 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1261;

architecture SYN_PLUTO_architecture208 of FD_1261 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2086 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2086);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture208;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1260 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1260;

architecture SYN_PLUTO_architecture209 of FD_1260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2087 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2087);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture209;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1259 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1259;

architecture SYN_PLUTO_architecture210 of FD_1259 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2088 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2088);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture210;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1258 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1258;

architecture SYN_PLUTO_architecture211 of FD_1258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2089 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2089);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture211;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1257 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1257;

architecture SYN_PLUTO_architecture212 of FD_1257 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2090 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2090);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture212;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1256 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1256;

architecture SYN_PLUTO_architecture213 of FD_1256 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2091 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2091);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture213;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1255 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1255;

architecture SYN_PLUTO_architecture214 of FD_1255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2092 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2092);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture214;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1254 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1254;

architecture SYN_PLUTO_architecture215 of FD_1254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2093 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2093);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture215;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1253 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1253;

architecture SYN_PLUTO_architecture216 of FD_1253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2094 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2094);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture216;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1252 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1252;

architecture SYN_PLUTO_architecture217 of FD_1252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2095 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2095);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture217;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1251 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1251;

architecture SYN_PLUTO_architecture218 of FD_1251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2096 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2096);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture218;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1250 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1250;

architecture SYN_PLUTO_architecture219 of FD_1250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2097 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2097);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture219;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1249 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1249;

architecture SYN_PLUTO_architecture220 of FD_1249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2098 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2098);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture220;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1248 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1248;

architecture SYN_PLUTO_architecture221 of FD_1248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2099 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2099);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture221;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1247 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1247;

architecture SYN_PLUTO_architecture222 of FD_1247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2100 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2100);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture222;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1246 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1246;

architecture SYN_PLUTO_architecture223 of FD_1246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2101 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2101);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture223;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1245 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1245;

architecture SYN_PLUTO_architecture224 of FD_1245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2102 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2102);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture224;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1244 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1244;

architecture SYN_PLUTO_architecture225 of FD_1244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2103 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2103);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture225;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1243 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1243;

architecture SYN_PLUTO_architecture226 of FD_1243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2104 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2104);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture226;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1242 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1242;

architecture SYN_PLUTO_architecture227 of FD_1242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2105 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2105);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture227;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1241 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1241;

architecture SYN_PLUTO_architecture228 of FD_1241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2106 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2106);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture228;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1240 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1240;

architecture SYN_PLUTO_architecture229 of FD_1240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2107 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2107);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture229;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1239 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1239;

architecture SYN_PLUTO_architecture230 of FD_1239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2108 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2108);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture230;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1238 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1238;

architecture SYN_PLUTO_architecture231 of FD_1238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2109 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2109);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture231;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1237 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1237;

architecture SYN_PLUTO_architecture232 of FD_1237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2110 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2110);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture232;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1236 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1236;

architecture SYN_PLUTO_architecture233 of FD_1236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2111 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2111);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture233;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1235 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1235;

architecture SYN_PLUTO_architecture234 of FD_1235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2112 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2112);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture234;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1234 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1234;

architecture SYN_PLUTO_architecture235 of FD_1234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2113 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2113);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture235;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1233 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1233;

architecture SYN_PLUTO_architecture236 of FD_1233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2114 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2114);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture236;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1232 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1232;

architecture SYN_PLUTO_architecture237 of FD_1232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2115 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2115);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture237;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1231 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1231;

architecture SYN_PLUTO_architecture238 of FD_1231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2116 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2116);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture238;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1230 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1230;

architecture SYN_PLUTO_architecture239 of FD_1230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2117 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2117);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture239;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1229 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1229;

architecture SYN_PLUTO_architecture240 of FD_1229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2118 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2118);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture240;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1228 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1228;

architecture SYN_PLUTO_architecture241 of FD_1228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2119 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2119);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture241;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1227 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1227;

architecture SYN_PLUTO_architecture242 of FD_1227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2120 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2120);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture242;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1226 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1226;

architecture SYN_PLUTO_architecture243 of FD_1226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2121 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2121);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture243;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1225 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1225;

architecture SYN_PLUTO_architecture244 of FD_1225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2122 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2122);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture244;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1224 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1224;

architecture SYN_PLUTO_architecture245 of FD_1224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2123 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2123);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture245;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1223 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1223;

architecture SYN_PLUTO_architecture246 of FD_1223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2124 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2124);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture246;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1222 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1222;

architecture SYN_PLUTO_architecture247 of FD_1222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2125 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2125);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture247;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1221 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1221;

architecture SYN_PLUTO_architecture248 of FD_1221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2126 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2126);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture248;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1220 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1220;

architecture SYN_PLUTO of FD_1220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2127 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2127);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1219 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1219;

architecture SYN_PLUTO_architecture of FD_1219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2128 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2128);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1218 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1218;

architecture SYN_PLUTO_architecture2 of FD_1218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2129 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2129);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1217 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1217;

architecture SYN_PLUTO_architecture3 of FD_1217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2130 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2130);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1216 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1216;

architecture SYN_PLUTO_architecture4 of FD_1216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2131 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2131);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1215 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1215;

architecture SYN_PLUTO_architecture5 of FD_1215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2132 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2132);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1214 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1214;

architecture SYN_PLUTO_architecture6 of FD_1214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2133 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2133);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1213 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1213;

architecture SYN_PLUTO_architecture7 of FD_1213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2134 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2134);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1212 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1212;

architecture SYN_PLUTO_architecture8 of FD_1212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2135 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2135);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1211 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1211;

architecture SYN_PLUTO_architecture9 of FD_1211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2136 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2136);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1210 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1210;

architecture SYN_PLUTO_architecture10 of FD_1210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2137 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2137);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1209 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1209;

architecture SYN_PLUTO_architecture11 of FD_1209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2138 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2138);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1208 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1208;

architecture SYN_PLUTO_architecture12 of FD_1208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2139 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2139);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1207 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1207;

architecture SYN_PLUTO_architecture13 of FD_1207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2140 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2140);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1206 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1206;

architecture SYN_PLUTO_architecture14 of FD_1206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2141 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2141);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1205 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1205;

architecture SYN_PLUTO_architecture15 of FD_1205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2142 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2142);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1204 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1204;

architecture SYN_PLUTO_architecture16 of FD_1204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2143 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2143);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1203 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1203;

architecture SYN_PLUTO_architecture17 of FD_1203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2144 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2144);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1202 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1202;

architecture SYN_PLUTO_architecture18 of FD_1202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2145 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2145);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1201 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1201;

architecture SYN_PLUTO_architecture19 of FD_1201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2146 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2146);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1200 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1200;

architecture SYN_PLUTO_architecture20 of FD_1200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2147 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2147);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1199 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1199;

architecture SYN_PLUTO_architecture21 of FD_1199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2148 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2148);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1198 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1198;

architecture SYN_PLUTO_architecture22 of FD_1198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2149 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2149);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1197 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1197;

architecture SYN_PLUTO_architecture23 of FD_1197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2150 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2150);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1196 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1196;

architecture SYN_PLUTO_architecture24 of FD_1196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2151 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2151);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1195 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1195;

architecture SYN_PLUTO_architecture25 of FD_1195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2152 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2152);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1194 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1194;

architecture SYN_PLUTO_architecture26 of FD_1194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2153 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2153);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1193 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1193;

architecture SYN_PLUTO_architecture27 of FD_1193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2154 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2154);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1192 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1192;

architecture SYN_PLUTO_architecture28 of FD_1192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2155 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2155);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1191 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1191;

architecture SYN_PLUTO_architecture29 of FD_1191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2156 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2156);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1190 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1190;

architecture SYN_PLUTO_architecture30 of FD_1190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2157 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2157);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1189 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1189;

architecture SYN_PLUTO_architecture31 of FD_1189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2158 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2158);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1188 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1188;

architecture SYN_PLUTO of FD_1188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2159 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2159);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1187 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1187;

architecture SYN_PLUTO_architecture of FD_1187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2160 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2160);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1186 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1186;

architecture SYN_PLUTO_architecture2 of FD_1186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2161 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2161);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1185 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1185;

architecture SYN_PLUTO_architecture3 of FD_1185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2162 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2162);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1184 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1184;

architecture SYN_PLUTO_architecture4 of FD_1184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2163 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2163);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1183 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1183;

architecture SYN_PLUTO_architecture5 of FD_1183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2164 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2164);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1182 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1182;

architecture SYN_PLUTO_architecture6 of FD_1182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2165 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2165);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1181 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1181;

architecture SYN_PLUTO_architecture7 of FD_1181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2166 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2166);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1180 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1180;

architecture SYN_PLUTO_architecture8 of FD_1180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2167 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2167);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1179 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1179;

architecture SYN_PLUTO_architecture9 of FD_1179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2168 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2168);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1178 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1178;

architecture SYN_PLUTO_architecture10 of FD_1178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2169 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2169);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1177 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1177;

architecture SYN_PLUTO_architecture11 of FD_1177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2170 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2170);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1176 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1176;

architecture SYN_PLUTO_architecture12 of FD_1176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2171 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2171);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1175 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1175;

architecture SYN_PLUTO_architecture13 of FD_1175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2172 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2172);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1174 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1174;

architecture SYN_PLUTO_architecture14 of FD_1174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2173 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2173);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1173 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1173;

architecture SYN_PLUTO_architecture15 of FD_1173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2174 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2174);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1172 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1172;

architecture SYN_PLUTO_architecture16 of FD_1172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2175 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2175);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1171 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1171;

architecture SYN_PLUTO_architecture17 of FD_1171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2176 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2176);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1170 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1170;

architecture SYN_PLUTO_architecture18 of FD_1170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2177 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2177);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1169 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1169;

architecture SYN_PLUTO_architecture19 of FD_1169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2178 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2178);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1168 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1168;

architecture SYN_PLUTO_architecture20 of FD_1168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2179 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2179);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1167 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1167;

architecture SYN_PLUTO_architecture21 of FD_1167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2180 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2180);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1166 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1166;

architecture SYN_PLUTO_architecture22 of FD_1166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2181 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2181);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1165 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1165;

architecture SYN_PLUTO_architecture23 of FD_1165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2182 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2182);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1164 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1164;

architecture SYN_PLUTO_architecture24 of FD_1164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2183 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2183);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1163 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1163;

architecture SYN_PLUTO_architecture25 of FD_1163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2184 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2184);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1162 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1162;

architecture SYN_PLUTO_architecture26 of FD_1162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2185 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2185);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1161 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1161;

architecture SYN_PLUTO_architecture27 of FD_1161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2186 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2186);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1160 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1160;

architecture SYN_PLUTO_architecture28 of FD_1160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2187 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2187);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1159 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1159;

architecture SYN_PLUTO_architecture29 of FD_1159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2188 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2188);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1158 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1158;

architecture SYN_PLUTO_architecture30 of FD_1158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2189 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2189);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1157 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1157;

architecture SYN_PLUTO_architecture31 of FD_1157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2190 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2190);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1156 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1156;

architecture SYN_PLUTO_architecture32 of FD_1156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2191 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2191);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1155 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1155;

architecture SYN_PLUTO_architecture33 of FD_1155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2192 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2192);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1154 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1154;

architecture SYN_PLUTO_architecture34 of FD_1154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2193 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2193);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1153 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1153;

architecture SYN_PLUTO_architecture35 of FD_1153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2194 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2194);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1152 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1152;

architecture SYN_PLUTO_architecture36 of FD_1152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2195 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2195);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1151 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1151;

architecture SYN_PLUTO_architecture37 of FD_1151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2196 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2196);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1150 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1150;

architecture SYN_PLUTO_architecture38 of FD_1150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2197 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2197);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1149 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1149;

architecture SYN_PLUTO_architecture39 of FD_1149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2198 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2198);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1148 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1148;

architecture SYN_PLUTO_architecture40 of FD_1148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2199 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2199);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1147 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1147;

architecture SYN_PLUTO_architecture41 of FD_1147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2200 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2200);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1146 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1146;

architecture SYN_PLUTO_architecture42 of FD_1146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2201 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2201);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1145 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1145;

architecture SYN_PLUTO_architecture43 of FD_1145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2202 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2202);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1144 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1144;

architecture SYN_PLUTO_architecture44 of FD_1144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2203 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2203);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1143 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1143;

architecture SYN_PLUTO_architecture45 of FD_1143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2204 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2204);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1142 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1142;

architecture SYN_PLUTO_architecture46 of FD_1142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2205 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2205);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1141 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1141;

architecture SYN_PLUTO_architecture47 of FD_1141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2206 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2206);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1140 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1140;

architecture SYN_PLUTO_architecture48 of FD_1140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2207 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2207);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1139 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1139;

architecture SYN_PLUTO_architecture49 of FD_1139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2208 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2208);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1138 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1138;

architecture SYN_PLUTO_architecture50 of FD_1138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2209 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2209);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1137 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1137;

architecture SYN_PLUTO_architecture51 of FD_1137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2210 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2210);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1136 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1136;

architecture SYN_PLUTO_architecture52 of FD_1136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2211 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2211);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1135 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1135;

architecture SYN_PLUTO_architecture53 of FD_1135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2212 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2212);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1134 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1134;

architecture SYN_PLUTO_architecture54 of FD_1134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2213 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2213);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1133 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1133;

architecture SYN_PLUTO_architecture55 of FD_1133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2214 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2214);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1132 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1132;

architecture SYN_PLUTO_architecture56 of FD_1132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2215 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2215);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1131 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1131;

architecture SYN_PLUTO_architecture57 of FD_1131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2216 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2216);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1130 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1130;

architecture SYN_PLUTO_architecture58 of FD_1130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2217 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2217);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1129 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1129;

architecture SYN_PLUTO_architecture59 of FD_1129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2218 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2218);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1128 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1128;

architecture SYN_PLUTO_architecture60 of FD_1128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2219 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2219);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1127 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1127;

architecture SYN_PLUTO_architecture61 of FD_1127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2220 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2220);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1126 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1126;

architecture SYN_PLUTO_architecture62 of FD_1126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2221 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2221);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1125 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1125;

architecture SYN_PLUTO_architecture63 of FD_1125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2222 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2222);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1124 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1124;

architecture SYN_PLUTO_architecture64 of FD_1124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2223 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2223);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1123 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1123;

architecture SYN_PLUTO_architecture65 of FD_1123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2224 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2224);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1122 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1122;

architecture SYN_PLUTO_architecture66 of FD_1122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2225 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2225);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1121 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1121;

architecture SYN_PLUTO_architecture67 of FD_1121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2226 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2226);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1120 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1120;

architecture SYN_PLUTO_architecture68 of FD_1120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2227 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2227);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1119 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1119;

architecture SYN_PLUTO_architecture69 of FD_1119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2228 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2228);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1118 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1118;

architecture SYN_PLUTO_architecture70 of FD_1118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2229 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2229);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1117 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1117;

architecture SYN_PLUTO_architecture71 of FD_1117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2230 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2230);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1116 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1116;

architecture SYN_PLUTO_architecture72 of FD_1116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2231 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2231);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1115 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1115;

architecture SYN_PLUTO_architecture73 of FD_1115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2232 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2232);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1114 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1114;

architecture SYN_PLUTO_architecture74 of FD_1114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2233 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2233);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1113 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1113;

architecture SYN_PLUTO_architecture75 of FD_1113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2234 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2234);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1112 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1112;

architecture SYN_PLUTO_architecture76 of FD_1112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2235 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2235);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1111 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1111;

architecture SYN_PLUTO_architecture77 of FD_1111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2236 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2236);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1110 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1110;

architecture SYN_PLUTO_architecture78 of FD_1110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2237 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2237);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1109 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1109;

architecture SYN_PLUTO_architecture79 of FD_1109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2238 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2238);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1108 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1108;

architecture SYN_PLUTO_architecture80 of FD_1108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2239 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2239);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1107 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1107;

architecture SYN_PLUTO_architecture81 of FD_1107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2240 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2240);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1106 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1106;

architecture SYN_PLUTO_architecture82 of FD_1106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2241 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2241);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1105 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1105;

architecture SYN_PLUTO_architecture83 of FD_1105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2242 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2242);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1104 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1104;

architecture SYN_PLUTO_architecture84 of FD_1104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2243 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2243);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1103 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1103;

architecture SYN_PLUTO_architecture85 of FD_1103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2244 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2244);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1102 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1102;

architecture SYN_PLUTO_architecture86 of FD_1102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2245 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2245);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1101 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1101;

architecture SYN_PLUTO_architecture87 of FD_1101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2246 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2246);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1100 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1100;

architecture SYN_PLUTO_architecture88 of FD_1100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2247 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2247);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1099 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1099;

architecture SYN_PLUTO_architecture89 of FD_1099 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2248 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2248);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1098 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1098;

architecture SYN_PLUTO_architecture90 of FD_1098 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2249 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2249);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1097 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1097;

architecture SYN_PLUTO_architecture91 of FD_1097 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2250 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2250);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1096 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1096;

architecture SYN_PLUTO_architecture92 of FD_1096 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2251 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2251);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1095 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1095;

architecture SYN_PLUTO_architecture93 of FD_1095 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2252 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2252);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1094 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1094;

architecture SYN_PLUTO_architecture94 of FD_1094 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2253 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2253);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1093 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1093;

architecture SYN_PLUTO_architecture95 of FD_1093 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2254 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2254);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1092 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1092;

architecture SYN_PLUTO_architecture96 of FD_1092 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2255 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2255);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1091 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1091;

architecture SYN_PLUTO_architecture97 of FD_1091 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2256 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2256);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1090 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1090;

architecture SYN_PLUTO_architecture98 of FD_1090 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2257 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2257);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1089 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1089;

architecture SYN_PLUTO_architecture99 of FD_1089 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2258 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2258);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1088 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1088;

architecture SYN_PLUTO_architecture100 of FD_1088 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2259 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2259);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1087 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1087;

architecture SYN_PLUTO_architecture101 of FD_1087 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2260 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2260);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1086 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1086;

architecture SYN_PLUTO_architecture102 of FD_1086 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2261 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2261);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1085 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1085;

architecture SYN_PLUTO_architecture103 of FD_1085 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2262 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2262);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1084 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1084;

architecture SYN_PLUTO_architecture104 of FD_1084 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2263 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2263);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1083 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1083;

architecture SYN_PLUTO_architecture105 of FD_1083 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2264 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2264);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1082 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1082;

architecture SYN_PLUTO_architecture106 of FD_1082 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2265 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2265);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1081 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1081;

architecture SYN_PLUTO_architecture107 of FD_1081 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2266 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2266);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1080 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1080;

architecture SYN_PLUTO_architecture108 of FD_1080 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2267 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2267);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1079 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1079;

architecture SYN_PLUTO_architecture109 of FD_1079 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2268 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2268);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1078 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1078;

architecture SYN_PLUTO_architecture110 of FD_1078 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2269 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2269);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1077 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1077;

architecture SYN_PLUTO_architecture111 of FD_1077 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2270 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2270);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1076 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1076;

architecture SYN_PLUTO_architecture112 of FD_1076 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2271 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2271);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1075 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1075;

architecture SYN_PLUTO_architecture113 of FD_1075 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2272 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2272);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1074 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1074;

architecture SYN_PLUTO_architecture114 of FD_1074 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2273 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2273);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1073 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1073;

architecture SYN_PLUTO_architecture115 of FD_1073 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2274 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2274);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1072 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1072;

architecture SYN_PLUTO_architecture116 of FD_1072 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2275 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2275);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1071 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1071;

architecture SYN_PLUTO_architecture117 of FD_1071 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2276 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2276);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1070 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1070;

architecture SYN_PLUTO_architecture118 of FD_1070 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2277 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2277);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1069 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1069;

architecture SYN_PLUTO_architecture119 of FD_1069 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2278 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2278);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1068 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1068;

architecture SYN_PLUTO_architecture120 of FD_1068 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2279 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2279);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1067 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1067;

architecture SYN_PLUTO_architecture121 of FD_1067 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2280 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2280);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1066 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1066;

architecture SYN_PLUTO_architecture122 of FD_1066 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2281 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2281);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1065 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1065;

architecture SYN_PLUTO_architecture123 of FD_1065 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2282 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2282);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1064 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1064;

architecture SYN_PLUTO_architecture124 of FD_1064 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2283 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2283);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1063 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1063;

architecture SYN_PLUTO_architecture125 of FD_1063 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2284 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2284);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1062 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1062;

architecture SYN_PLUTO_architecture126 of FD_1062 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2285 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2285);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1061 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1061;

architecture SYN_PLUTO_architecture127 of FD_1061 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2286 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2286);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1060 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1060;

architecture SYN_PLUTO_architecture128 of FD_1060 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2287 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2287);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1059 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1059;

architecture SYN_PLUTO_architecture129 of FD_1059 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2288 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2288);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1058 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1058;

architecture SYN_PLUTO_architecture130 of FD_1058 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2289 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2289);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1057 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1057;

architecture SYN_PLUTO_architecture131 of FD_1057 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2290 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2290);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1056 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1056;

architecture SYN_PLUTO_architecture132 of FD_1056 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2291 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2291);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1055 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1055;

architecture SYN_PLUTO_architecture133 of FD_1055 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2292 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2292);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1054 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1054;

architecture SYN_PLUTO_architecture134 of FD_1054 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2293 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2293);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1053 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1053;

architecture SYN_PLUTO_architecture135 of FD_1053 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2294 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2294);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1052 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1052;

architecture SYN_PLUTO_architecture136 of FD_1052 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2295 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2295);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1051 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1051;

architecture SYN_PLUTO_architecture137 of FD_1051 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2296 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2296);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1050 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1050;

architecture SYN_PLUTO_architecture138 of FD_1050 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2297 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2297);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1049 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1049;

architecture SYN_PLUTO_architecture139 of FD_1049 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2298 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2298);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1048 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1048;

architecture SYN_PLUTO_architecture140 of FD_1048 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2299 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2299);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1047 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1047;

architecture SYN_PLUTO_architecture141 of FD_1047 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2300 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2300);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1046 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1046;

architecture SYN_PLUTO_architecture142 of FD_1046 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2301 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2301);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1045 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1045;

architecture SYN_PLUTO_architecture143 of FD_1045 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2302 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2302);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture143;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1044 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1044;

architecture SYN_PLUTO_architecture144 of FD_1044 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2303 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2303);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture144;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1043 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1043;

architecture SYN_PLUTO_architecture145 of FD_1043 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2304 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2304);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture145;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1042 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1042;

architecture SYN_PLUTO_architecture146 of FD_1042 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2305 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2305);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture146;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1041 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1041;

architecture SYN_PLUTO_architecture147 of FD_1041 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2306 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2306);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture147;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1040 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1040;

architecture SYN_PLUTO_architecture148 of FD_1040 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2307 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2307);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture148;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1039 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1039;

architecture SYN_PLUTO_architecture149 of FD_1039 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2308 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2308);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture149;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1038 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1038;

architecture SYN_PLUTO_architecture150 of FD_1038 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2309 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2309);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture150;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1037 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1037;

architecture SYN_PLUTO_architecture151 of FD_1037 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2310 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2310);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture151;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1036 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1036;

architecture SYN_PLUTO_architecture152 of FD_1036 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2311 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2311);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture152;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1035 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1035;

architecture SYN_PLUTO_architecture153 of FD_1035 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2312 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2312);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture153;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1034 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1034;

architecture SYN_PLUTO_architecture154 of FD_1034 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2313 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2313);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture154;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1033 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1033;

architecture SYN_PLUTO_architecture155 of FD_1033 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2314 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2314);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture155;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1032 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1032;

architecture SYN_PLUTO_architecture156 of FD_1032 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2315 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2315);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture156;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1031 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1031;

architecture SYN_PLUTO_architecture157 of FD_1031 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2316 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2316);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture157;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1030 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1030;

architecture SYN_PLUTO_architecture158 of FD_1030 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2317 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2317);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture158;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1029 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1029;

architecture SYN_PLUTO_architecture159 of FD_1029 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2318 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2318);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture159;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1028 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1028;

architecture SYN_PLUTO_architecture160 of FD_1028 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2319 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2319);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture160;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1027 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1027;

architecture SYN_PLUTO_architecture161 of FD_1027 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2320 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2320);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture161;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1026 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1026;

architecture SYN_PLUTO_architecture162 of FD_1026 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2321 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2321);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture162;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1025 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1025;

architecture SYN_PLUTO_architecture163 of FD_1025 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2322 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2322);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture163;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1024 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1024;

architecture SYN_PLUTO_architecture164 of FD_1024 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2323 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2323);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture164;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1023 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1023;

architecture SYN_PLUTO_architecture165 of FD_1023 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2324 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2324);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture165;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1022 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1022;

architecture SYN_PLUTO_architecture166 of FD_1022 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2325 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2325);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture166;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1021 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1021;

architecture SYN_PLUTO_architecture167 of FD_1021 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2326 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2326);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture167;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1020 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1020;

architecture SYN_PLUTO_architecture168 of FD_1020 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2327 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2327);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture168;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1019 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1019;

architecture SYN_PLUTO_architecture169 of FD_1019 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2328 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2328);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture169;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1018 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1018;

architecture SYN_PLUTO_architecture170 of FD_1018 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2329 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2329);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture170;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1017 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1017;

architecture SYN_PLUTO_architecture171 of FD_1017 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2330 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2330);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture171;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1016 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1016;

architecture SYN_PLUTO_architecture172 of FD_1016 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2331 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2331);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture172;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1015 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1015;

architecture SYN_PLUTO_architecture173 of FD_1015 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2332 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2332);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture173;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1014 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1014;

architecture SYN_PLUTO_architecture174 of FD_1014 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2333 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2333);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture174;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1013 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1013;

architecture SYN_PLUTO_architecture175 of FD_1013 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2334 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2334);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture175;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1012 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1012;

architecture SYN_PLUTO_architecture176 of FD_1012 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2335 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2335);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture176;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1011 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1011;

architecture SYN_PLUTO_architecture177 of FD_1011 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2336 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2336);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture177;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1010 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1010;

architecture SYN_PLUTO_architecture178 of FD_1010 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2337 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2337);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture178;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1009 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1009;

architecture SYN_PLUTO_architecture179 of FD_1009 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2338 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2338);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture179;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1008 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1008;

architecture SYN_PLUTO_architecture180 of FD_1008 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2339 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2339);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture180;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1007 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1007;

architecture SYN_PLUTO_architecture181 of FD_1007 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2340 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2340);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture181;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1006 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1006;

architecture SYN_PLUTO_architecture182 of FD_1006 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2341 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2341);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture182;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1005 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1005;

architecture SYN_PLUTO_architecture183 of FD_1005 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2342 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2342);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture183;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1004 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1004;

architecture SYN_PLUTO_architecture184 of FD_1004 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2343 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2343);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture184;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1003 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1003;

architecture SYN_PLUTO_architecture185 of FD_1003 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2344 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2344);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture185;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1002 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1002;

architecture SYN_PLUTO_architecture186 of FD_1002 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2345 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2345);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture186;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1001 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1001;

architecture SYN_PLUTO_architecture187 of FD_1001 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2346 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2346);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture187;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1000 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1000;

architecture SYN_PLUTO_architecture188 of FD_1000 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2347 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2347);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture188;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_999 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_999;

architecture SYN_PLUTO_architecture189 of FD_999 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2348 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2348);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture189;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_998 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_998;

architecture SYN_PLUTO_architecture190 of FD_998 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2349 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2349);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture190;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_997 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_997;

architecture SYN_PLUTO_architecture191 of FD_997 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2350 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2350);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture191;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_996 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_996;

architecture SYN_PLUTO_architecture192 of FD_996 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2351 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2351);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture192;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_995 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_995;

architecture SYN_PLUTO_architecture193 of FD_995 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2352 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2352);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture193;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_994 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_994;

architecture SYN_PLUTO_architecture194 of FD_994 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2353 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2353);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture194;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_993 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_993;

architecture SYN_PLUTO_architecture195 of FD_993 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2354 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2354);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture195;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_992 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_992;

architecture SYN_PLUTO_architecture196 of FD_992 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2355 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2355);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture196;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_991 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_991;

architecture SYN_PLUTO_architecture197 of FD_991 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2356 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2356);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture197;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_990 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_990;

architecture SYN_PLUTO_architecture198 of FD_990 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2357 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2357);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture198;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_989 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_989;

architecture SYN_PLUTO_architecture199 of FD_989 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2358 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2358);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture199;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_988 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_988;

architecture SYN_PLUTO_architecture200 of FD_988 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2359 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2359);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture200;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_987 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_987;

architecture SYN_PLUTO_architecture201 of FD_987 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2360 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2360);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture201;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_986 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_986;

architecture SYN_PLUTO_architecture202 of FD_986 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2361 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2361);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture202;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_985 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_985;

architecture SYN_PLUTO_architecture203 of FD_985 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2362 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2362);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture203;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_984 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_984;

architecture SYN_PLUTO_architecture204 of FD_984 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2363 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2363);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture204;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_983 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_983;

architecture SYN_PLUTO_architecture205 of FD_983 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2364 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2364);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture205;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_982 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_982;

architecture SYN_PLUTO_architecture206 of FD_982 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2365 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2365);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture206;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_981 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_981;

architecture SYN_PLUTO_architecture207 of FD_981 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2366 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2366);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture207;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_980 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_980;

architecture SYN_PLUTO_architecture208 of FD_980 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2367 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2367);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture208;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_979 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_979;

architecture SYN_PLUTO_architecture209 of FD_979 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2368 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2368);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture209;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_978 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_978;

architecture SYN_PLUTO_architecture210 of FD_978 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2369 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2369);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture210;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_977 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_977;

architecture SYN_PLUTO_architecture211 of FD_977 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2370 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2370);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture211;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_976 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_976;

architecture SYN_PLUTO_architecture212 of FD_976 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2371 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2371);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture212;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_975 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_975;

architecture SYN_PLUTO_architecture213 of FD_975 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2372 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2372);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture213;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_974 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_974;

architecture SYN_PLUTO_architecture214 of FD_974 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2373 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2373);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture214;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_973 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_973;

architecture SYN_PLUTO_architecture215 of FD_973 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2374 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2374);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture215;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_972 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_972;

architecture SYN_PLUTO_architecture216 of FD_972 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2375 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2375);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture216;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_971 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_971;

architecture SYN_PLUTO_architecture217 of FD_971 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2376 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2376);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture217;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_970 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_970;

architecture SYN_PLUTO_architecture218 of FD_970 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2377 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2377);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture218;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_969 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_969;

architecture SYN_PLUTO_architecture219 of FD_969 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2378 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2378);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture219;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_968 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_968;

architecture SYN_PLUTO_architecture220 of FD_968 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2379 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2379);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture220;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_967 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_967;

architecture SYN_PLUTO_architecture221 of FD_967 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2380 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2380);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture221;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_966 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_966;

architecture SYN_PLUTO_architecture222 of FD_966 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2381 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2381);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture222;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_965 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_965;

architecture SYN_PLUTO_architecture223 of FD_965 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2382 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2382);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture223;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_964 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_964;

architecture SYN_PLUTO_architecture224 of FD_964 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2383 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2383);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture224;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_963 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_963;

architecture SYN_PLUTO_architecture225 of FD_963 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2384 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2384);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture225;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_962 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_962;

architecture SYN_PLUTO_architecture226 of FD_962 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2385 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2385);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture226;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_961 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_961;

architecture SYN_PLUTO_architecture227 of FD_961 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2386 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2386);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture227;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_960 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_960;

architecture SYN_PLUTO_architecture228 of FD_960 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2387 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2387);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture228;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_959 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_959;

architecture SYN_PLUTO_architecture229 of FD_959 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2388 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2388);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture229;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_958 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_958;

architecture SYN_PLUTO_architecture230 of FD_958 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2389 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2389);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture230;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_957 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_957;

architecture SYN_PLUTO_architecture231 of FD_957 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2390 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2390);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture231;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_956 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_956;

architecture SYN_PLUTO_architecture232 of FD_956 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2391 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2391);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture232;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_955 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_955;

architecture SYN_PLUTO_architecture233 of FD_955 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2392 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2392);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture233;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_954 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_954;

architecture SYN_PLUTO_architecture234 of FD_954 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2393 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2393);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture234;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_953 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_953;

architecture SYN_PLUTO_architecture235 of FD_953 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2394 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2394);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture235;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_952 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_952;

architecture SYN_PLUTO_architecture236 of FD_952 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2395 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2395);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture236;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_951 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_951;

architecture SYN_PLUTO_architecture237 of FD_951 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2396 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2396);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture237;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_950 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_950;

architecture SYN_PLUTO_architecture238 of FD_950 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2397 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2397);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture238;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_949 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_949;

architecture SYN_PLUTO_architecture239 of FD_949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2398 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2398);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture239;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_948 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_948;

architecture SYN_PLUTO_architecture240 of FD_948 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2399 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2399);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture240;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_947 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_947;

architecture SYN_PLUTO_architecture241 of FD_947 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2400 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2400);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture241;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_946 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_946;

architecture SYN_PLUTO_architecture242 of FD_946 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2401 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2401);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture242;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_945 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_945;

architecture SYN_PLUTO_architecture243 of FD_945 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2402 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2402);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture243;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_944 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_944;

architecture SYN_PLUTO_architecture244 of FD_944 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2403 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2403);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture244;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_943 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_943;

architecture SYN_PLUTO_architecture245 of FD_943 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2404 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2404);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture245;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_942 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_942;

architecture SYN_PLUTO_architecture246 of FD_942 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2405 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2405);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture246;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_941 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_941;

architecture SYN_PLUTO_architecture247 of FD_941 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2406 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2406);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture247;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_940 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_940;

architecture SYN_PLUTO_architecture248 of FD_940 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2407 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2407);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture248;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_939 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_939;

architecture SYN_PLUTO of FD_939 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2408 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2408);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_938 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_938;

architecture SYN_PLUTO_architecture of FD_938 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2409 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2409);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_937 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_937;

architecture SYN_PLUTO_architecture2 of FD_937 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2410 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2410);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_936 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_936;

architecture SYN_PLUTO_architecture3 of FD_936 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2411 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2411);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_935 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_935;

architecture SYN_PLUTO_architecture4 of FD_935 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2412 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2412);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_934 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_934;

architecture SYN_PLUTO_architecture5 of FD_934 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2413 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2413);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_933 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_933;

architecture SYN_PLUTO_architecture6 of FD_933 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2414 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2414);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_932 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_932;

architecture SYN_PLUTO_architecture7 of FD_932 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2415 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2415);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_931 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_931;

architecture SYN_PLUTO_architecture8 of FD_931 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2416 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2416);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_930 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_930;

architecture SYN_PLUTO_architecture9 of FD_930 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2417 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2417);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_929 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_929;

architecture SYN_PLUTO_architecture10 of FD_929 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2418 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2418);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_928 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_928;

architecture SYN_PLUTO_architecture11 of FD_928 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2419 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2419);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_927 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_927;

architecture SYN_PLUTO_architecture12 of FD_927 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2420 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2420);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_926 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_926;

architecture SYN_PLUTO_architecture13 of FD_926 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2421 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2421);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_925 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_925;

architecture SYN_PLUTO_architecture14 of FD_925 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2422 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2422);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_924 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_924;

architecture SYN_PLUTO_architecture15 of FD_924 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2423 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2423);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_923 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_923;

architecture SYN_PLUTO_architecture16 of FD_923 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2424 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2424);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_922 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_922;

architecture SYN_PLUTO_architecture17 of FD_922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2425 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2425);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_921 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_921;

architecture SYN_PLUTO_architecture18 of FD_921 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2426 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2426);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_920 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_920;

architecture SYN_PLUTO_architecture19 of FD_920 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2427 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2427);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_919 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_919;

architecture SYN_PLUTO_architecture20 of FD_919 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2428 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2428);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_918 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_918;

architecture SYN_PLUTO_architecture21 of FD_918 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2429 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2429);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_917 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_917;

architecture SYN_PLUTO_architecture22 of FD_917 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2430 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2430);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_916 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_916;

architecture SYN_PLUTO_architecture23 of FD_916 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2431 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2431);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_915 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_915;

architecture SYN_PLUTO_architecture24 of FD_915 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2432 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2432);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_914 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_914;

architecture SYN_PLUTO_architecture25 of FD_914 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2433 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2433);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_913 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_913;

architecture SYN_PLUTO_architecture26 of FD_913 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2434 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2434);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_912 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_912;

architecture SYN_PLUTO_architecture27 of FD_912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2435 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2435);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_911 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_911;

architecture SYN_PLUTO_architecture28 of FD_911 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2436 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2436);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_910 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_910;

architecture SYN_PLUTO_architecture29 of FD_910 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2437 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2437);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_909 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_909;

architecture SYN_PLUTO_architecture30 of FD_909 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2438 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2438);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_908 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_908;

architecture SYN_PLUTO_architecture31 of FD_908 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2439 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2439);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_907 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_907;

architecture SYN_PLUTO of FD_907 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2440 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2440);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_906 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_906;

architecture SYN_PLUTO_architecture of FD_906 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2441 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2441);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_905 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_905;

architecture SYN_PLUTO_architecture2 of FD_905 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2442 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2442);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_904 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_904;

architecture SYN_PLUTO_architecture3 of FD_904 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2443 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2443);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_903 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_903;

architecture SYN_PLUTO_architecture4 of FD_903 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2444 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2444);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_902 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_902;

architecture SYN_PLUTO_architecture5 of FD_902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2445 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2445);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_901 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_901;

architecture SYN_PLUTO_architecture6 of FD_901 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2446 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2446);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_900 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_900;

architecture SYN_PLUTO_architecture7 of FD_900 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2447 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2447);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_899 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_899;

architecture SYN_PLUTO_architecture8 of FD_899 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2448 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2448);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_898 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_898;

architecture SYN_PLUTO_architecture9 of FD_898 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2449 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2449);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_897 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_897;

architecture SYN_PLUTO_architecture10 of FD_897 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2450 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2450);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_896 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_896;

architecture SYN_PLUTO_architecture11 of FD_896 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2451 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2451);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_895 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_895;

architecture SYN_PLUTO_architecture12 of FD_895 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2452 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2452);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_894 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_894;

architecture SYN_PLUTO_architecture13 of FD_894 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2453 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2453);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_893 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_893;

architecture SYN_PLUTO_architecture14 of FD_893 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2454 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2454);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_892 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_892;

architecture SYN_PLUTO_architecture15 of FD_892 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2455 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2455);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_891 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_891;

architecture SYN_PLUTO_architecture16 of FD_891 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2456 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2456);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_890 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_890;

architecture SYN_PLUTO_architecture17 of FD_890 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2457 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2457);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_889 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_889;

architecture SYN_PLUTO_architecture18 of FD_889 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2458 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2458);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_888 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_888;

architecture SYN_PLUTO_architecture19 of FD_888 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2459 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2459);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_887 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_887;

architecture SYN_PLUTO_architecture20 of FD_887 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2460 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2460);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_886 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_886;

architecture SYN_PLUTO_architecture21 of FD_886 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2461 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2461);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_885 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_885;

architecture SYN_PLUTO_architecture22 of FD_885 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2462 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2462);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_884 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_884;

architecture SYN_PLUTO_architecture23 of FD_884 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2463 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2463);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_883 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_883;

architecture SYN_PLUTO_architecture24 of FD_883 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2464 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2464);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_882 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_882;

architecture SYN_PLUTO_architecture25 of FD_882 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2465 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2465);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_881 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_881;

architecture SYN_PLUTO_architecture26 of FD_881 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2466 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2466);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_880 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_880;

architecture SYN_PLUTO_architecture27 of FD_880 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2467 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2467);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_879 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_879;

architecture SYN_PLUTO_architecture28 of FD_879 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2468 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2468);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_878 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_878;

architecture SYN_PLUTO_architecture29 of FD_878 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2469 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2469);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_877 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_877;

architecture SYN_PLUTO_architecture30 of FD_877 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2470 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2470);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_876 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_876;

architecture SYN_PLUTO_architecture31 of FD_876 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2471 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2471);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_875 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_875;

architecture SYN_PLUTO_architecture32 of FD_875 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2472 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2472);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_874 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_874;

architecture SYN_PLUTO_architecture33 of FD_874 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2473 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2473);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_873 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_873;

architecture SYN_PLUTO_architecture34 of FD_873 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2474 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2474);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_872 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_872;

architecture SYN_PLUTO_architecture35 of FD_872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2475 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2475);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_871 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_871;

architecture SYN_PLUTO_architecture36 of FD_871 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2476 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2476);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_870 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_870;

architecture SYN_PLUTO_architecture37 of FD_870 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2477 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2477);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_869 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_869;

architecture SYN_PLUTO_architecture38 of FD_869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2478 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2478);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_868 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_868;

architecture SYN_PLUTO_architecture39 of FD_868 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2479 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2479);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_867 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_867;

architecture SYN_PLUTO_architecture40 of FD_867 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2480 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2480);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_866 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_866;

architecture SYN_PLUTO_architecture41 of FD_866 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2481 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2481);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_865 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_865;

architecture SYN_PLUTO_architecture42 of FD_865 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2482 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2482);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_864 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_864;

architecture SYN_PLUTO_architecture43 of FD_864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2483 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2483);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_863 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_863;

architecture SYN_PLUTO_architecture44 of FD_863 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2484 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2484);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_862 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_862;

architecture SYN_PLUTO_architecture45 of FD_862 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2485 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2485);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_861 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_861;

architecture SYN_PLUTO_architecture46 of FD_861 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2486 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2486);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_860 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_860;

architecture SYN_PLUTO_architecture47 of FD_860 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2487 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2487);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_859 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_859;

architecture SYN_PLUTO_architecture48 of FD_859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2488 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2488);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_858 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_858;

architecture SYN_PLUTO_architecture49 of FD_858 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2489 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2489);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_857 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_857;

architecture SYN_PLUTO_architecture50 of FD_857 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2490 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2490);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_856 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_856;

architecture SYN_PLUTO_architecture51 of FD_856 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2491 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2491);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_855 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_855;

architecture SYN_PLUTO_architecture52 of FD_855 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2492 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2492);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_854 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_854;

architecture SYN_PLUTO_architecture53 of FD_854 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2493 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2493);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_853 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_853;

architecture SYN_PLUTO_architecture54 of FD_853 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2494 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2494);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_852 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_852;

architecture SYN_PLUTO_architecture55 of FD_852 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2495 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2495);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_851 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_851;

architecture SYN_PLUTO_architecture56 of FD_851 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2496 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2496);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_850 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_850;

architecture SYN_PLUTO_architecture57 of FD_850 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2497 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2497);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_849 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_849;

architecture SYN_PLUTO_architecture58 of FD_849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2498 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2498);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_848 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_848;

architecture SYN_PLUTO_architecture59 of FD_848 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2499 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2499);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_847 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_847;

architecture SYN_PLUTO_architecture60 of FD_847 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2500 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2500);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_846 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_846;

architecture SYN_PLUTO_architecture61 of FD_846 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2501 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2501);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_845 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_845;

architecture SYN_PLUTO_architecture62 of FD_845 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2502 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2502);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_844 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_844;

architecture SYN_PLUTO_architecture63 of FD_844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2503 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2503);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_843 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_843;

architecture SYN_PLUTO_architecture64 of FD_843 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2504 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2504);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_842 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_842;

architecture SYN_PLUTO_architecture65 of FD_842 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2505 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2505);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_841 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_841;

architecture SYN_PLUTO_architecture66 of FD_841 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2506 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2506);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_840 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_840;

architecture SYN_PLUTO_architecture67 of FD_840 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2507 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2507);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_839 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_839;

architecture SYN_PLUTO_architecture68 of FD_839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2508 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2508);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_838 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_838;

architecture SYN_PLUTO_architecture69 of FD_838 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2509 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2509);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_837 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_837;

architecture SYN_PLUTO_architecture70 of FD_837 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2510 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2510);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_836 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_836;

architecture SYN_PLUTO_architecture71 of FD_836 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2511 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2511);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_835 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_835;

architecture SYN_PLUTO_architecture72 of FD_835 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2512 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2512);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_834 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_834;

architecture SYN_PLUTO_architecture73 of FD_834 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2513 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2513);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_833 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_833;

architecture SYN_PLUTO_architecture74 of FD_833 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2514 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2514);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_832 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_832;

architecture SYN_PLUTO_architecture75 of FD_832 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2515 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2515);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_831 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_831;

architecture SYN_PLUTO_architecture76 of FD_831 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2516 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2516);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_830 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_830;

architecture SYN_PLUTO_architecture77 of FD_830 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2517 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2517);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_829 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_829;

architecture SYN_PLUTO_architecture78 of FD_829 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2518 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2518);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_828 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_828;

architecture SYN_PLUTO_architecture79 of FD_828 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2519 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2519);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_827 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_827;

architecture SYN_PLUTO_architecture80 of FD_827 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2520 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2520);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_826 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_826;

architecture SYN_PLUTO_architecture81 of FD_826 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2521 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2521);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_825 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_825;

architecture SYN_PLUTO_architecture82 of FD_825 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2522 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2522);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_824 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_824;

architecture SYN_PLUTO_architecture83 of FD_824 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2523 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2523);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_823 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_823;

architecture SYN_PLUTO_architecture84 of FD_823 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2524 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2524);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_822 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_822;

architecture SYN_PLUTO_architecture85 of FD_822 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2525 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2525);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_821 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_821;

architecture SYN_PLUTO_architecture86 of FD_821 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2526 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2526);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_820 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_820;

architecture SYN_PLUTO_architecture87 of FD_820 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2527 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2527);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_819 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_819;

architecture SYN_PLUTO_architecture88 of FD_819 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2528 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2528);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_818 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_818;

architecture SYN_PLUTO_architecture89 of FD_818 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2529 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2529);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_817 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_817;

architecture SYN_PLUTO_architecture90 of FD_817 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2530 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2530);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_816 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_816;

architecture SYN_PLUTO_architecture91 of FD_816 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2531 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2531);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_815 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_815;

architecture SYN_PLUTO_architecture92 of FD_815 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2532 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2532);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_814 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_814;

architecture SYN_PLUTO_architecture93 of FD_814 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2533 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2533);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_813 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_813;

architecture SYN_PLUTO_architecture94 of FD_813 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2534 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2534);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_812 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_812;

architecture SYN_PLUTO_architecture95 of FD_812 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2535 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2535);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_811 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_811;

architecture SYN_PLUTO_architecture96 of FD_811 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2536 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2536);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_810 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_810;

architecture SYN_PLUTO_architecture97 of FD_810 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2537 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2537);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_809 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_809;

architecture SYN_PLUTO_architecture98 of FD_809 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2538 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2538);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_808 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_808;

architecture SYN_PLUTO_architecture99 of FD_808 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2539 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2539);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_807 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_807;

architecture SYN_PLUTO_architecture100 of FD_807 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2540 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2540);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_806 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_806;

architecture SYN_PLUTO_architecture101 of FD_806 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2541 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2541);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_805 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_805;

architecture SYN_PLUTO_architecture102 of FD_805 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2542 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2542);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_804 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_804;

architecture SYN_PLUTO_architecture103 of FD_804 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2543 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2543);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_803 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_803;

architecture SYN_PLUTO_architecture104 of FD_803 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2544 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2544);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_802 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_802;

architecture SYN_PLUTO_architecture105 of FD_802 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2545 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2545);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_801 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_801;

architecture SYN_PLUTO_architecture106 of FD_801 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2546 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2546);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_800 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_800;

architecture SYN_PLUTO_architecture107 of FD_800 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2547 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2547);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_799 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_799;

architecture SYN_PLUTO_architecture108 of FD_799 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2548 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2548);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_798 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_798;

architecture SYN_PLUTO_architecture109 of FD_798 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2549 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2549);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_797 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_797;

architecture SYN_PLUTO_architecture110 of FD_797 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2550 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2550);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_796 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_796;

architecture SYN_PLUTO_architecture111 of FD_796 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2551 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2551);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_795 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_795;

architecture SYN_PLUTO_architecture112 of FD_795 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2552 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2552);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_794 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_794;

architecture SYN_PLUTO_architecture113 of FD_794 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2553 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2553);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_793 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_793;

architecture SYN_PLUTO_architecture114 of FD_793 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2554 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2554);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_792 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_792;

architecture SYN_PLUTO_architecture115 of FD_792 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2555 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2555);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_791 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_791;

architecture SYN_PLUTO_architecture116 of FD_791 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2556 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2556);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_790 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_790;

architecture SYN_PLUTO_architecture117 of FD_790 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2557 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2557);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_789 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_789;

architecture SYN_PLUTO_architecture118 of FD_789 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2558 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2558);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_788 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_788;

architecture SYN_PLUTO_architecture119 of FD_788 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2559 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2559);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_787 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_787;

architecture SYN_PLUTO_architecture120 of FD_787 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2560 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2560);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_786 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_786;

architecture SYN_PLUTO_architecture121 of FD_786 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2561 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2561);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_785 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_785;

architecture SYN_PLUTO_architecture122 of FD_785 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2562 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2562);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_784 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_784;

architecture SYN_PLUTO_architecture123 of FD_784 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2563 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2563);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_783 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_783;

architecture SYN_PLUTO_architecture124 of FD_783 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2564 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2564);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_782 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_782;

architecture SYN_PLUTO_architecture125 of FD_782 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2565 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2565);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_781 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_781;

architecture SYN_PLUTO_architecture126 of FD_781 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2566 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2566);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_780 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_780;

architecture SYN_PLUTO_architecture127 of FD_780 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2567 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2567);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_779 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_779;

architecture SYN_PLUTO_architecture128 of FD_779 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2568 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2568);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_778 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_778;

architecture SYN_PLUTO_architecture129 of FD_778 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2569 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2569);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_777 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_777;

architecture SYN_PLUTO_architecture130 of FD_777 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2570 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2570);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_776 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_776;

architecture SYN_PLUTO_architecture131 of FD_776 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2571 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2571);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_775 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_775;

architecture SYN_PLUTO_architecture132 of FD_775 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2572 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2572);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_774 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_774;

architecture SYN_PLUTO_architecture133 of FD_774 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2573 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2573);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_773 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_773;

architecture SYN_PLUTO_architecture134 of FD_773 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2574 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2574);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_772 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_772;

architecture SYN_PLUTO_architecture135 of FD_772 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2575 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2575);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_771 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_771;

architecture SYN_PLUTO_architecture136 of FD_771 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2576 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2576);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_770 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_770;

architecture SYN_PLUTO_architecture137 of FD_770 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2577 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2577);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_769 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_769;

architecture SYN_PLUTO_architecture138 of FD_769 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2578 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2578);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_768 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_768;

architecture SYN_PLUTO_architecture139 of FD_768 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2579 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2579);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_767 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_767;

architecture SYN_PLUTO_architecture140 of FD_767 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2580 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2580);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_766 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_766;

architecture SYN_PLUTO_architecture141 of FD_766 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2581 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2581);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_765 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_765;

architecture SYN_PLUTO_architecture142 of FD_765 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2582 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2582);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_764 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_764;

architecture SYN_PLUTO_architecture143 of FD_764 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2583 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2583);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture143;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_763 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_763;

architecture SYN_PLUTO_architecture144 of FD_763 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2584 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2584);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture144;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_762 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_762;

architecture SYN_PLUTO_architecture145 of FD_762 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2585 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2585);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture145;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_761 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_761;

architecture SYN_PLUTO_architecture146 of FD_761 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2586 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2586);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture146;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_760 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_760;

architecture SYN_PLUTO_architecture147 of FD_760 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2587 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2587);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture147;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_759 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_759;

architecture SYN_PLUTO_architecture148 of FD_759 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2588 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2588);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture148;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_758 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_758;

architecture SYN_PLUTO_architecture149 of FD_758 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2589 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2589);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture149;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_757 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_757;

architecture SYN_PLUTO_architecture150 of FD_757 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2590 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2590);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture150;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_756 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_756;

architecture SYN_PLUTO_architecture151 of FD_756 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2591 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2591);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture151;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_755 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_755;

architecture SYN_PLUTO_architecture152 of FD_755 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2592 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2592);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture152;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_754 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_754;

architecture SYN_PLUTO_architecture153 of FD_754 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2593 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2593);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture153;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_753 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_753;

architecture SYN_PLUTO_architecture154 of FD_753 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2594 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2594);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture154;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_752 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_752;

architecture SYN_PLUTO_architecture155 of FD_752 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2595 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2595);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture155;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_751 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_751;

architecture SYN_PLUTO_architecture156 of FD_751 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2596 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2596);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture156;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_750 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_750;

architecture SYN_PLUTO_architecture157 of FD_750 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2597 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2597);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture157;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_749 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_749;

architecture SYN_PLUTO_architecture158 of FD_749 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2598 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2598);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture158;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_748 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_748;

architecture SYN_PLUTO_architecture159 of FD_748 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2599 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2599);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture159;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_747 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_747;

architecture SYN_PLUTO_architecture160 of FD_747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2600 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2600);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture160;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_746 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_746;

architecture SYN_PLUTO_architecture161 of FD_746 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2601 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2601);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture161;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_745 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_745;

architecture SYN_PLUTO_architecture162 of FD_745 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2602 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2602);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture162;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_744 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_744;

architecture SYN_PLUTO_architecture163 of FD_744 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2603 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2603);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture163;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_743 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_743;

architecture SYN_PLUTO_architecture164 of FD_743 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2604 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2604);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture164;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_742 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_742;

architecture SYN_PLUTO_architecture165 of FD_742 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2605 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2605);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture165;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_741 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_741;

architecture SYN_PLUTO_architecture166 of FD_741 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2606 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2606);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture166;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_740 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_740;

architecture SYN_PLUTO_architecture167 of FD_740 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2607 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2607);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture167;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_739 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_739;

architecture SYN_PLUTO_architecture168 of FD_739 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2608 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2608);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture168;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_738 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_738;

architecture SYN_PLUTO_architecture169 of FD_738 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2609 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2609);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture169;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_737 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_737;

architecture SYN_PLUTO_architecture170 of FD_737 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2610 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2610);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture170;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_736 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_736;

architecture SYN_PLUTO_architecture171 of FD_736 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2611 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2611);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture171;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_735 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_735;

architecture SYN_PLUTO_architecture172 of FD_735 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2612 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2612);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture172;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_734 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_734;

architecture SYN_PLUTO_architecture173 of FD_734 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2613 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2613);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture173;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_733 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_733;

architecture SYN_PLUTO_architecture174 of FD_733 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2614 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2614);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture174;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_732 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_732;

architecture SYN_PLUTO_architecture175 of FD_732 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2615 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2615);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture175;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_731 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_731;

architecture SYN_PLUTO_architecture176 of FD_731 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2616 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2616);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture176;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_730 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_730;

architecture SYN_PLUTO_architecture177 of FD_730 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2617 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2617);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture177;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_729 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_729;

architecture SYN_PLUTO_architecture178 of FD_729 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2618 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2618);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture178;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_728 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_728;

architecture SYN_PLUTO_architecture179 of FD_728 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2619 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2619);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture179;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_727 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_727;

architecture SYN_PLUTO_architecture180 of FD_727 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2620 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2620);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture180;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_726 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_726;

architecture SYN_PLUTO_architecture181 of FD_726 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2621 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2621);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture181;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_725 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_725;

architecture SYN_PLUTO_architecture182 of FD_725 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2622 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2622);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture182;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_724 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_724;

architecture SYN_PLUTO_architecture183 of FD_724 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2623 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2623);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture183;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_723 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_723;

architecture SYN_PLUTO_architecture184 of FD_723 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2624 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2624);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture184;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_722 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_722;

architecture SYN_PLUTO_architecture185 of FD_722 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2625 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2625);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture185;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_721 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_721;

architecture SYN_PLUTO_architecture186 of FD_721 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2626 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2626);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture186;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_720 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_720;

architecture SYN_PLUTO_architecture187 of FD_720 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2627 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2627);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture187;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_719 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_719;

architecture SYN_PLUTO_architecture188 of FD_719 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2628 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2628);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture188;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_718 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_718;

architecture SYN_PLUTO_architecture189 of FD_718 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2629 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2629);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture189;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_717 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_717;

architecture SYN_PLUTO_architecture190 of FD_717 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2630 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2630);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture190;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_716 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_716;

architecture SYN_PLUTO_architecture191 of FD_716 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2631 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2631);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture191;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_715 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_715;

architecture SYN_PLUTO_architecture192 of FD_715 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2632 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2632);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture192;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_714 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_714;

architecture SYN_PLUTO_architecture193 of FD_714 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2633 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2633);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture193;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_713 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_713;

architecture SYN_PLUTO_architecture194 of FD_713 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2634 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2634);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture194;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_712 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_712;

architecture SYN_PLUTO_architecture195 of FD_712 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2635 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2635);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture195;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_711 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_711;

architecture SYN_PLUTO_architecture196 of FD_711 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2636 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2636);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture196;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_710 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_710;

architecture SYN_PLUTO_architecture197 of FD_710 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2637 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2637);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture197;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_709 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_709;

architecture SYN_PLUTO_architecture198 of FD_709 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2638 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2638);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture198;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_708 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_708;

architecture SYN_PLUTO_architecture199 of FD_708 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2639 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2639);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture199;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_707 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_707;

architecture SYN_PLUTO_architecture200 of FD_707 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2640 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2640);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture200;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_706 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_706;

architecture SYN_PLUTO_architecture201 of FD_706 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2641 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2641);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture201;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_705 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_705;

architecture SYN_PLUTO_architecture202 of FD_705 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2642 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2642);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture202;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_704 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_704;

architecture SYN_PLUTO_architecture203 of FD_704 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2643 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2643);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture203;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_703 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_703;

architecture SYN_PLUTO_architecture204 of FD_703 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2644 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2644);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture204;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_702 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_702;

architecture SYN_PLUTO_architecture205 of FD_702 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2645 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2645);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture205;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_701 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_701;

architecture SYN_PLUTO_architecture206 of FD_701 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2646 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2646);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture206;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_700 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_700;

architecture SYN_PLUTO_architecture207 of FD_700 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2647 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2647);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture207;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_699 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_699;

architecture SYN_PLUTO_architecture208 of FD_699 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2648 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2648);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture208;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_698 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_698;

architecture SYN_PLUTO_architecture209 of FD_698 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2649 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2649);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture209;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_697 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_697;

architecture SYN_PLUTO_architecture210 of FD_697 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2650 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2650);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture210;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_696 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_696;

architecture SYN_PLUTO_architecture211 of FD_696 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2651 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2651);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture211;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_695 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_695;

architecture SYN_PLUTO_architecture212 of FD_695 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2652 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2652);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture212;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_694 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_694;

architecture SYN_PLUTO_architecture213 of FD_694 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2653 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2653);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture213;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_693 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_693;

architecture SYN_PLUTO_architecture214 of FD_693 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2654 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2654);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture214;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_692 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_692;

architecture SYN_PLUTO_architecture215 of FD_692 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2655 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2655);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture215;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_691 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_691;

architecture SYN_PLUTO_architecture216 of FD_691 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2656 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2656);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture216;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_690 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_690;

architecture SYN_PLUTO_architecture217 of FD_690 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2657 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2657);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture217;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_689 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_689;

architecture SYN_PLUTO_architecture218 of FD_689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2658 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2658);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture218;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_688 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_688;

architecture SYN_PLUTO_architecture219 of FD_688 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2659 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2659);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture219;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_687 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_687;

architecture SYN_PLUTO_architecture220 of FD_687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2660 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2660);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture220;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_686 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_686;

architecture SYN_PLUTO_architecture221 of FD_686 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2661 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2661);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture221;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_685 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_685;

architecture SYN_PLUTO_architecture222 of FD_685 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2662 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2662);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture222;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_684 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_684;

architecture SYN_PLUTO_architecture223 of FD_684 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2663 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2663);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture223;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_683 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_683;

architecture SYN_PLUTO_architecture224 of FD_683 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2664 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2664);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture224;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_682 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_682;

architecture SYN_PLUTO_architecture225 of FD_682 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2665 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2665);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture225;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_681 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_681;

architecture SYN_PLUTO_architecture226 of FD_681 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2666 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2666);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture226;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_680 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_680;

architecture SYN_PLUTO_architecture227 of FD_680 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2667 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2667);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture227;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_679 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_679;

architecture SYN_PLUTO_architecture228 of FD_679 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2668 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2668);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture228;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_678 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_678;

architecture SYN_PLUTO_architecture229 of FD_678 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2669 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2669);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture229;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_677 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_677;

architecture SYN_PLUTO_architecture230 of FD_677 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2670 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2670);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture230;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_676 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_676;

architecture SYN_PLUTO_architecture231 of FD_676 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2671 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2671);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture231;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_675 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_675;

architecture SYN_PLUTO_architecture232 of FD_675 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2672 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2672);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture232;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_674 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_674;

architecture SYN_PLUTO_architecture233 of FD_674 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2673 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2673);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture233;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_673 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_673;

architecture SYN_PLUTO_architecture234 of FD_673 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2674 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2674);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture234;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_672 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_672;

architecture SYN_PLUTO_architecture235 of FD_672 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2675 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2675);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture235;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_671 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_671;

architecture SYN_PLUTO_architecture236 of FD_671 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2676 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2676);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture236;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_670 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_670;

architecture SYN_PLUTO_architecture237 of FD_670 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2677 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2677);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture237;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_669 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_669;

architecture SYN_PLUTO_architecture238 of FD_669 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2678 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2678);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture238;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_668 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_668;

architecture SYN_PLUTO_architecture239 of FD_668 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2679 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2679);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture239;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_667 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_667;

architecture SYN_PLUTO_architecture240 of FD_667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2680 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2680);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture240;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_666 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_666;

architecture SYN_PLUTO_architecture241 of FD_666 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2681 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2681);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture241;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_665 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_665;

architecture SYN_PLUTO_architecture242 of FD_665 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2682 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2682);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture242;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_664 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_664;

architecture SYN_PLUTO_architecture243 of FD_664 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2683 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2683);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture243;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_663 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_663;

architecture SYN_PLUTO_architecture244 of FD_663 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2684 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2684);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture244;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_662 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_662;

architecture SYN_PLUTO_architecture245 of FD_662 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2685 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2685);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture245;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_661 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_661;

architecture SYN_PLUTO_architecture246 of FD_661 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2686 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2686);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture246;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_660 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_660;

architecture SYN_PLUTO_architecture247 of FD_660 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2687 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2687);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture247;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_659 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_659;

architecture SYN_PLUTO_architecture248 of FD_659 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2688 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2688);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture248;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_658 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_658;

architecture SYN_PLUTO of FD_658 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2689 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2689);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_657 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_657;

architecture SYN_PLUTO_architecture of FD_657 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2690 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2690);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_656 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_656;

architecture SYN_PLUTO_architecture2 of FD_656 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2691 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2691);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_655 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_655;

architecture SYN_PLUTO_architecture3 of FD_655 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2692 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2692);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_654 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_654;

architecture SYN_PLUTO_architecture4 of FD_654 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2693 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2693);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_653 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_653;

architecture SYN_PLUTO_architecture5 of FD_653 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2694 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2694);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_652 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_652;

architecture SYN_PLUTO_architecture6 of FD_652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2695 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2695);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_651 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_651;

architecture SYN_PLUTO_architecture7 of FD_651 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2696 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2696);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_650 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_650;

architecture SYN_PLUTO_architecture8 of FD_650 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2697 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2697);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_649 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_649;

architecture SYN_PLUTO_architecture9 of FD_649 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2698 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2698);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_648 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_648;

architecture SYN_PLUTO_architecture10 of FD_648 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2699 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2699);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_647 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_647;

architecture SYN_PLUTO_architecture11 of FD_647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2700 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2700);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_646 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_646;

architecture SYN_PLUTO_architecture12 of FD_646 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2701 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2701);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_645 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_645;

architecture SYN_PLUTO_architecture13 of FD_645 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2702 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2702);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_644 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_644;

architecture SYN_PLUTO_architecture14 of FD_644 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2703 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2703);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_643 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_643;

architecture SYN_PLUTO_architecture15 of FD_643 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2704 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2704);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_642 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_642;

architecture SYN_PLUTO_architecture16 of FD_642 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2705 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2705);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_641 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_641;

architecture SYN_PLUTO_architecture17 of FD_641 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2706 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2706);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_640 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_640;

architecture SYN_PLUTO_architecture18 of FD_640 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2707 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2707);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_639 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_639;

architecture SYN_PLUTO_architecture19 of FD_639 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2708 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2708);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_638 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_638;

architecture SYN_PLUTO_architecture20 of FD_638 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2709 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2709);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_637 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_637;

architecture SYN_PLUTO_architecture21 of FD_637 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2710 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2710);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_636 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_636;

architecture SYN_PLUTO_architecture22 of FD_636 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2711 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2711);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_635 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_635;

architecture SYN_PLUTO_architecture23 of FD_635 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2712 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2712);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_634 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_634;

architecture SYN_PLUTO_architecture24 of FD_634 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2713 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2713);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_633 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_633;

architecture SYN_PLUTO_architecture25 of FD_633 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2714 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2714);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_632 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_632;

architecture SYN_PLUTO_architecture26 of FD_632 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2715 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2715);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_631 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_631;

architecture SYN_PLUTO_architecture27 of FD_631 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2716 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2716);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_630 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_630;

architecture SYN_PLUTO_architecture28 of FD_630 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2717 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2717);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_629 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_629;

architecture SYN_PLUTO_architecture29 of FD_629 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2718 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2718);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_628 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_628;

architecture SYN_PLUTO_architecture30 of FD_628 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2719 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2719);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_627 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_627;

architecture SYN_PLUTO_architecture31 of FD_627 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2720 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2720);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_626 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_626;

architecture SYN_PLUTO of FD_626 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2721 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2721);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_625 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_625;

architecture SYN_PLUTO_architecture of FD_625 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2722 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2722);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_624 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_624;

architecture SYN_PLUTO_architecture2 of FD_624 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2723 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2723);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_623 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_623;

architecture SYN_PLUTO_architecture3 of FD_623 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2724 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2724);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_622 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_622;

architecture SYN_PLUTO_architecture4 of FD_622 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2725 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2725);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_621 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_621;

architecture SYN_PLUTO_architecture5 of FD_621 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2726 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2726);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_620 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_620;

architecture SYN_PLUTO_architecture6 of FD_620 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2727 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2727);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_619 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_619;

architecture SYN_PLUTO_architecture7 of FD_619 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2728 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2728);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_618 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_618;

architecture SYN_PLUTO_architecture8 of FD_618 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2729 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2729);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_617 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_617;

architecture SYN_PLUTO_architecture9 of FD_617 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2730 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2730);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_616 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_616;

architecture SYN_PLUTO_architecture10 of FD_616 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2731 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2731);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_615 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_615;

architecture SYN_PLUTO_architecture11 of FD_615 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2732 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2732);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_614 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_614;

architecture SYN_PLUTO_architecture12 of FD_614 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2733 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2733);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_613 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_613;

architecture SYN_PLUTO_architecture13 of FD_613 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2734 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2734);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_612 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_612;

architecture SYN_PLUTO_architecture14 of FD_612 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2735 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2735);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_611 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_611;

architecture SYN_PLUTO_architecture15 of FD_611 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2736 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2736);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_610 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_610;

architecture SYN_PLUTO_architecture16 of FD_610 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2737 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2737);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_609 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_609;

architecture SYN_PLUTO_architecture17 of FD_609 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2738 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2738);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_608 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_608;

architecture SYN_PLUTO_architecture18 of FD_608 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2739 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2739);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_607 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_607;

architecture SYN_PLUTO_architecture19 of FD_607 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2740 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2740);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_606 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_606;

architecture SYN_PLUTO_architecture20 of FD_606 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2741 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2741);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_605 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_605;

architecture SYN_PLUTO_architecture21 of FD_605 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2742 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2742);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_604 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_604;

architecture SYN_PLUTO_architecture22 of FD_604 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2743 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2743);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_603 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_603;

architecture SYN_PLUTO_architecture23 of FD_603 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2744 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2744);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_602 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_602;

architecture SYN_PLUTO_architecture24 of FD_602 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2745 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2745);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_601 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_601;

architecture SYN_PLUTO_architecture25 of FD_601 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2746 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2746);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_600 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_600;

architecture SYN_PLUTO_architecture26 of FD_600 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2747 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2747);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_599 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_599;

architecture SYN_PLUTO_architecture27 of FD_599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2748 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2748);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_598 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_598;

architecture SYN_PLUTO_architecture28 of FD_598 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2749 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2749);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_597 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_597;

architecture SYN_PLUTO_architecture29 of FD_597 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2750 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2750);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_596 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_596;

architecture SYN_PLUTO_architecture30 of FD_596 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2751 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2751);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_595 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_595;

architecture SYN_PLUTO_architecture31 of FD_595 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2752 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2752);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_594 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_594;

architecture SYN_PLUTO_architecture32 of FD_594 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2753 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2753);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_593 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_593;

architecture SYN_PLUTO_architecture33 of FD_593 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2754 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2754);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_592 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_592;

architecture SYN_PLUTO_architecture34 of FD_592 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2755 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2755);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_591 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_591;

architecture SYN_PLUTO_architecture35 of FD_591 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2756 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2756);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_590 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_590;

architecture SYN_PLUTO_architecture36 of FD_590 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2757 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2757);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_589 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_589;

architecture SYN_PLUTO_architecture37 of FD_589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2758 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2758);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_588 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_588;

architecture SYN_PLUTO_architecture38 of FD_588 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2759 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2759);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_587 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_587;

architecture SYN_PLUTO_architecture39 of FD_587 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2760 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2760);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_586 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_586;

architecture SYN_PLUTO_architecture40 of FD_586 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2761 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2761);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_585 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_585;

architecture SYN_PLUTO_architecture41 of FD_585 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2762 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2762);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_584 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_584;

architecture SYN_PLUTO_architecture42 of FD_584 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2763 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2763);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_583 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_583;

architecture SYN_PLUTO_architecture43 of FD_583 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2764 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2764);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_582 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_582;

architecture SYN_PLUTO_architecture44 of FD_582 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2765 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2765);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_581 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_581;

architecture SYN_PLUTO_architecture45 of FD_581 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2766 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2766);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_580 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_580;

architecture SYN_PLUTO_architecture46 of FD_580 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2767 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2767);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_579 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_579;

architecture SYN_PLUTO_architecture47 of FD_579 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2768 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2768);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_578 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_578;

architecture SYN_PLUTO_architecture48 of FD_578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2769 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2769);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_577 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_577;

architecture SYN_PLUTO_architecture49 of FD_577 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2770 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2770);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_576 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_576;

architecture SYN_PLUTO_architecture50 of FD_576 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2771 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2771);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_575 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_575;

architecture SYN_PLUTO_architecture51 of FD_575 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2772 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2772);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_574 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_574;

architecture SYN_PLUTO_architecture52 of FD_574 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2773 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2773);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_573 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_573;

architecture SYN_PLUTO_architecture53 of FD_573 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2774 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2774);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_572 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_572;

architecture SYN_PLUTO_architecture54 of FD_572 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2775 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2775);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_571 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_571;

architecture SYN_PLUTO_architecture55 of FD_571 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2776 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2776);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_570 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_570;

architecture SYN_PLUTO_architecture56 of FD_570 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2777 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2777);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_569 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_569;

architecture SYN_PLUTO_architecture57 of FD_569 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2778 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2778);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_568 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_568;

architecture SYN_PLUTO_architecture58 of FD_568 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2779 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2779);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_567 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_567;

architecture SYN_PLUTO_architecture59 of FD_567 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2780 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2780);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_566 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_566;

architecture SYN_PLUTO_architecture60 of FD_566 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2781 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2781);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_565 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_565;

architecture SYN_PLUTO_architecture61 of FD_565 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2782 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2782);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_564 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_564;

architecture SYN_PLUTO_architecture62 of FD_564 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2783 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2783);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_563 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_563;

architecture SYN_PLUTO_architecture63 of FD_563 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2784 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2784);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_562 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_562;

architecture SYN_PLUTO_architecture64 of FD_562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2785 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2785);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_561 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_561;

architecture SYN_PLUTO_architecture65 of FD_561 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2786 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2786);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_560 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_560;

architecture SYN_PLUTO_architecture66 of FD_560 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2787 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2787);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_559 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_559;

architecture SYN_PLUTO_architecture67 of FD_559 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2788 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2788);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_558 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_558;

architecture SYN_PLUTO_architecture68 of FD_558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2789 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2789);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_557 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_557;

architecture SYN_PLUTO_architecture69 of FD_557 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2790 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2790);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_556 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_556;

architecture SYN_PLUTO_architecture70 of FD_556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2791 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2791);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_555 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_555;

architecture SYN_PLUTO_architecture71 of FD_555 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2792 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2792);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_554 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_554;

architecture SYN_PLUTO_architecture72 of FD_554 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2793 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2793);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_553 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_553;

architecture SYN_PLUTO_architecture73 of FD_553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2794 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2794);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_552 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_552;

architecture SYN_PLUTO_architecture74 of FD_552 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2795 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2795);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_551 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_551;

architecture SYN_PLUTO_architecture75 of FD_551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2796 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2796);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_550 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_550;

architecture SYN_PLUTO_architecture76 of FD_550 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2797 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2797);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_549 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_549;

architecture SYN_PLUTO_architecture77 of FD_549 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2798 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2798);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_548 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_548;

architecture SYN_PLUTO_architecture78 of FD_548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2799 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2799);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_547 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_547;

architecture SYN_PLUTO_architecture79 of FD_547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2800 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2800);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_546 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_546;

architecture SYN_PLUTO_architecture80 of FD_546 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2801 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2801);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_545 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_545;

architecture SYN_PLUTO_architecture81 of FD_545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2802 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2802);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_544 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_544;

architecture SYN_PLUTO_architecture82 of FD_544 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2803 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2803);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_543 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_543;

architecture SYN_PLUTO_architecture83 of FD_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2804 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2804);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_542 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_542;

architecture SYN_PLUTO_architecture84 of FD_542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2805 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2805);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_541 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_541;

architecture SYN_PLUTO_architecture85 of FD_541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2806 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2806);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_540 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_540;

architecture SYN_PLUTO_architecture86 of FD_540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2807 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2807);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_539 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_539;

architecture SYN_PLUTO_architecture87 of FD_539 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2808 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2808);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_538 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_538;

architecture SYN_PLUTO_architecture88 of FD_538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2809 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2809);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_537 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_537;

architecture SYN_PLUTO_architecture89 of FD_537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2810 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2810);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_536 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_536;

architecture SYN_PLUTO_architecture90 of FD_536 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2811 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2811);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_535 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_535;

architecture SYN_PLUTO_architecture91 of FD_535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2812 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2812);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_534 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_534;

architecture SYN_PLUTO_architecture92 of FD_534 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2813 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2813);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_533 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_533;

architecture SYN_PLUTO_architecture93 of FD_533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2814 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2814);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_532 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_532;

architecture SYN_PLUTO_architecture94 of FD_532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2815 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2815);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_531 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_531;

architecture SYN_PLUTO_architecture95 of FD_531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2816 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2816);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_530 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_530;

architecture SYN_PLUTO_architecture96 of FD_530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2817 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2817);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_529 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_529;

architecture SYN_PLUTO_architecture97 of FD_529 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2818 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2818);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_528 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_528;

architecture SYN_PLUTO_architecture98 of FD_528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2819 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2819);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_527 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_527;

architecture SYN_PLUTO_architecture99 of FD_527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2820 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2820);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_526 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_526;

architecture SYN_PLUTO_architecture100 of FD_526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2821 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2821);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_525 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_525;

architecture SYN_PLUTO_architecture101 of FD_525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2822 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2822);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_524 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_524;

architecture SYN_PLUTO_architecture102 of FD_524 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2823 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2823);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_523 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_523;

architecture SYN_PLUTO_architecture103 of FD_523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2824 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2824);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_522 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_522;

architecture SYN_PLUTO_architecture104 of FD_522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2825 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2825);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_521 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_521;

architecture SYN_PLUTO_architecture105 of FD_521 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2826 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2826);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_520 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_520;

architecture SYN_PLUTO_architecture106 of FD_520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2827 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2827);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_519 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_519;

architecture SYN_PLUTO_architecture107 of FD_519 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2828 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2828);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_518 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_518;

architecture SYN_PLUTO_architecture108 of FD_518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2829 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2829);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_517 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_517;

architecture SYN_PLUTO_architecture109 of FD_517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2830 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2830);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_516 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_516;

architecture SYN_PLUTO_architecture110 of FD_516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2831 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2831);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_515 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_515;

architecture SYN_PLUTO_architecture111 of FD_515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2832 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2832);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_514 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_514;

architecture SYN_PLUTO_architecture112 of FD_514 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2833 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2833);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_513 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_513;

architecture SYN_PLUTO_architecture113 of FD_513 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2834 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2834);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_512 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_512;

architecture SYN_PLUTO_architecture114 of FD_512 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2835 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2835);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_511 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_511;

architecture SYN_PLUTO_architecture115 of FD_511 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2836 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2836);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_510 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_510;

architecture SYN_PLUTO_architecture116 of FD_510 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2837 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2837);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_509 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_509;

architecture SYN_PLUTO_architecture117 of FD_509 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2838 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2838);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_508 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_508;

architecture SYN_PLUTO_architecture118 of FD_508 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2839 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2839);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_507 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_507;

architecture SYN_PLUTO_architecture119 of FD_507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2840 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2840);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_506 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_506;

architecture SYN_PLUTO_architecture120 of FD_506 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2841 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2841);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_505 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_505;

architecture SYN_PLUTO_architecture121 of FD_505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2842 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2842);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_504 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_504;

architecture SYN_PLUTO_architecture122 of FD_504 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2843 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2843);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_503 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_503;

architecture SYN_PLUTO_architecture123 of FD_503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2844 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2844);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_502 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_502;

architecture SYN_PLUTO_architecture124 of FD_502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2845 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2845);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_501 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_501;

architecture SYN_PLUTO_architecture125 of FD_501 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2846 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2846);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_500 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_500;

architecture SYN_PLUTO_architecture126 of FD_500 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2847 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2847);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_499 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_499;

architecture SYN_PLUTO_architecture127 of FD_499 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2848 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2848);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_498 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_498;

architecture SYN_PLUTO_architecture128 of FD_498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2849 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2849);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_497 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_497;

architecture SYN_PLUTO_architecture129 of FD_497 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2850 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2850);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_496 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_496;

architecture SYN_PLUTO_architecture130 of FD_496 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2851 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2851);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_495 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_495;

architecture SYN_PLUTO_architecture131 of FD_495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2852 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2852);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_494 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_494;

architecture SYN_PLUTO_architecture132 of FD_494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2853 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2853);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_493 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_493;

architecture SYN_PLUTO_architecture133 of FD_493 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2854 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2854);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_492 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_492;

architecture SYN_PLUTO_architecture134 of FD_492 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2855 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2855);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_491 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_491;

architecture SYN_PLUTO_architecture135 of FD_491 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2856 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2856);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_490 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_490;

architecture SYN_PLUTO_architecture136 of FD_490 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2857 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2857);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_489 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_489;

architecture SYN_PLUTO_architecture137 of FD_489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2858 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2858);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_488 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_488;

architecture SYN_PLUTO_architecture138 of FD_488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2859 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2859);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_487 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_487;

architecture SYN_PLUTO_architecture139 of FD_487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2860 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2860);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_486 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_486;

architecture SYN_PLUTO_architecture140 of FD_486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2861 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2861);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_485 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_485;

architecture SYN_PLUTO_architecture141 of FD_485 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2862 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2862);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_484 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_484;

architecture SYN_PLUTO_architecture142 of FD_484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2863 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2863);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_483 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_483;

architecture SYN_PLUTO_architecture143 of FD_483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2864 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2864);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture143;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_482 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_482;

architecture SYN_PLUTO_architecture144 of FD_482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2865 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2865);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture144;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_481 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_481;

architecture SYN_PLUTO_architecture145 of FD_481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2866 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2866);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture145;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_480 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_480;

architecture SYN_PLUTO_architecture146 of FD_480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2867 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2867);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture146;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_479 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_479;

architecture SYN_PLUTO_architecture147 of FD_479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2868 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2868);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture147;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_478 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_478;

architecture SYN_PLUTO_architecture148 of FD_478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2869 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2869);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture148;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_477 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_477;

architecture SYN_PLUTO_architecture149 of FD_477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2870 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2870);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture149;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_476 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_476;

architecture SYN_PLUTO_architecture150 of FD_476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2871 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2871);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture150;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_475 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_475;

architecture SYN_PLUTO_architecture151 of FD_475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2872 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2872);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture151;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_474 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_474;

architecture SYN_PLUTO_architecture152 of FD_474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2873 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2873);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture152;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_473 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_473;

architecture SYN_PLUTO_architecture153 of FD_473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2874 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2874);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture153;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_472 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_472;

architecture SYN_PLUTO_architecture154 of FD_472 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2875 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2875);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture154;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_471 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_471;

architecture SYN_PLUTO_architecture155 of FD_471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2876 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2876);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture155;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_470 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_470;

architecture SYN_PLUTO_architecture156 of FD_470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2877 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2877);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture156;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_469 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_469;

architecture SYN_PLUTO_architecture157 of FD_469 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2878 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2878);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture157;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_468 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_468;

architecture SYN_PLUTO_architecture158 of FD_468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2879 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2879);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture158;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_467 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_467;

architecture SYN_PLUTO_architecture159 of FD_467 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2880 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2880);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture159;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_466 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_466;

architecture SYN_PLUTO_architecture160 of FD_466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2881 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2881);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture160;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_465 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_465;

architecture SYN_PLUTO_architecture161 of FD_465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2882 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2882);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture161;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_464 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_464;

architecture SYN_PLUTO_architecture162 of FD_464 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2883 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2883);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture162;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_463 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_463;

architecture SYN_PLUTO_architecture163 of FD_463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2884 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2884);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture163;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_462 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_462;

architecture SYN_PLUTO_architecture164 of FD_462 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2885 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2885);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture164;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_461 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_461;

architecture SYN_PLUTO_architecture165 of FD_461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2886 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2886);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture165;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_460 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_460;

architecture SYN_PLUTO_architecture166 of FD_460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2887 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2887);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture166;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_459 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_459;

architecture SYN_PLUTO_architecture167 of FD_459 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2888 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2888);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture167;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_458 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_458;

architecture SYN_PLUTO_architecture168 of FD_458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2889 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2889);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture168;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_457 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_457;

architecture SYN_PLUTO_architecture169 of FD_457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2890 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2890);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture169;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_456 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_456;

architecture SYN_PLUTO_architecture170 of FD_456 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2891 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2891);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture170;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_455 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_455;

architecture SYN_PLUTO_architecture171 of FD_455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2892 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2892);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture171;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_454 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_454;

architecture SYN_PLUTO_architecture172 of FD_454 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2893 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2893);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture172;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_453 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_453;

architecture SYN_PLUTO_architecture173 of FD_453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2894 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2894);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture173;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_452 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_452;

architecture SYN_PLUTO_architecture174 of FD_452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2895 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2895);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture174;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_451 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_451;

architecture SYN_PLUTO_architecture175 of FD_451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2896 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2896);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture175;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_450 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_450;

architecture SYN_PLUTO_architecture176 of FD_450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2897 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2897);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture176;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_449 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_449;

architecture SYN_PLUTO_architecture177 of FD_449 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2898 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2898);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture177;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_448 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_448;

architecture SYN_PLUTO_architecture178 of FD_448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2899 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2899);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture178;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_447 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_447;

architecture SYN_PLUTO_architecture179 of FD_447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2900 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2900);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture179;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_446 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_446;

architecture SYN_PLUTO_architecture180 of FD_446 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2901 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2901);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture180;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_445 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_445;

architecture SYN_PLUTO_architecture181 of FD_445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2902 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2902);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture181;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_444 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_444;

architecture SYN_PLUTO_architecture182 of FD_444 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2903 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2903);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture182;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_443 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_443;

architecture SYN_PLUTO_architecture183 of FD_443 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2904 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2904);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture183;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_442 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_442;

architecture SYN_PLUTO_architecture184 of FD_442 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2905 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2905);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture184;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_441 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_441;

architecture SYN_PLUTO_architecture185 of FD_441 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2906 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2906);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture185;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_440 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_440;

architecture SYN_PLUTO_architecture186 of FD_440 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2907 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2907);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture186;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_439 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_439;

architecture SYN_PLUTO_architecture187 of FD_439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2908 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2908);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture187;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_438 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_438;

architecture SYN_PLUTO_architecture188 of FD_438 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2909 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2909);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture188;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_437 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_437;

architecture SYN_PLUTO_architecture189 of FD_437 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2910 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2910);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture189;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_436 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_436;

architecture SYN_PLUTO_architecture190 of FD_436 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2911 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2911);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture190;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_435 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_435;

architecture SYN_PLUTO_architecture191 of FD_435 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2912 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2912);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture191;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_434 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_434;

architecture SYN_PLUTO_architecture192 of FD_434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2913 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2913);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture192;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_433 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_433;

architecture SYN_PLUTO_architecture193 of FD_433 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2914 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2914);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture193;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_432 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_432;

architecture SYN_PLUTO_architecture194 of FD_432 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2915 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2915);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture194;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_431 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_431;

architecture SYN_PLUTO_architecture195 of FD_431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2916 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2916);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture195;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_430 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_430;

architecture SYN_PLUTO_architecture196 of FD_430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2917 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2917);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture196;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_429 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_429;

architecture SYN_PLUTO_architecture197 of FD_429 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2918 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2918);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture197;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_428 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_428;

architecture SYN_PLUTO_architecture198 of FD_428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2919 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2919);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture198;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_427 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_427;

architecture SYN_PLUTO_architecture199 of FD_427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2920 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2920);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture199;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_426 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_426;

architecture SYN_PLUTO_architecture200 of FD_426 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2921 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2921);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture200;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_425 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_425;

architecture SYN_PLUTO_architecture201 of FD_425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2922 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2922);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture201;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_424 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_424;

architecture SYN_PLUTO_architecture202 of FD_424 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2923 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2923);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture202;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_423 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_423;

architecture SYN_PLUTO_architecture203 of FD_423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2924 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2924);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture203;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_422 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_422;

architecture SYN_PLUTO_architecture204 of FD_422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2925 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2925);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture204;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_421 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_421;

architecture SYN_PLUTO_architecture205 of FD_421 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2926 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2926);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture205;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_420 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_420;

architecture SYN_PLUTO_architecture206 of FD_420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2927 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2927);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture206;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_419 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_419;

architecture SYN_PLUTO_architecture207 of FD_419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2928 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2928);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture207;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_418 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_418;

architecture SYN_PLUTO_architecture208 of FD_418 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2929 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2929);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture208;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_417 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_417;

architecture SYN_PLUTO_architecture209 of FD_417 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2930 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2930);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture209;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_416 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_416;

architecture SYN_PLUTO_architecture210 of FD_416 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2931 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2931);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture210;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_415 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_415;

architecture SYN_PLUTO_architecture211 of FD_415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2932 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2932);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture211;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_414 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_414;

architecture SYN_PLUTO_architecture212 of FD_414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2933 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2933);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture212;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_413 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_413;

architecture SYN_PLUTO_architecture213 of FD_413 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2934 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2934);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture213;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_412 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_412;

architecture SYN_PLUTO_architecture214 of FD_412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2935 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2935);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture214;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_411 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_411;

architecture SYN_PLUTO_architecture215 of FD_411 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2936 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2936);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture215;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_410 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_410;

architecture SYN_PLUTO_architecture216 of FD_410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2937 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2937);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture216;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_409 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_409;

architecture SYN_PLUTO_architecture217 of FD_409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2938 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2938);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture217;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_408 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_408;

architecture SYN_PLUTO_architecture218 of FD_408 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2939 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2939);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture218;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_407 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_407;

architecture SYN_PLUTO_architecture219 of FD_407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2940 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2940);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture219;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_406 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_406;

architecture SYN_PLUTO_architecture220 of FD_406 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2941 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2941);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture220;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_405 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_405;

architecture SYN_PLUTO_architecture221 of FD_405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2942 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2942);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture221;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_404 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_404;

architecture SYN_PLUTO_architecture222 of FD_404 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2943 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2943);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture222;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_403 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_403;

architecture SYN_PLUTO_architecture223 of FD_403 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2944 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2944);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture223;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_402 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_402;

architecture SYN_PLUTO_architecture224 of FD_402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2945 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2945);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture224;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_401 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_401;

architecture SYN_PLUTO_architecture225 of FD_401 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2946 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2946);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture225;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_400 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_400;

architecture SYN_PLUTO_architecture226 of FD_400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2947 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2947);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture226;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_399 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_399;

architecture SYN_PLUTO_architecture227 of FD_399 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2948 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2948);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture227;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_398 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_398;

architecture SYN_PLUTO_architecture228 of FD_398 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2949 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2949);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture228;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_397 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_397;

architecture SYN_PLUTO_architecture229 of FD_397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2950 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2950);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture229;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_396 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_396;

architecture SYN_PLUTO_architecture230 of FD_396 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2951 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2951);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture230;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_395 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_395;

architecture SYN_PLUTO_architecture231 of FD_395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2952 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2952);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture231;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_394 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_394;

architecture SYN_PLUTO_architecture232 of FD_394 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2953 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2953);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture232;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_393 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_393;

architecture SYN_PLUTO_architecture233 of FD_393 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2954 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2954);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture233;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_392 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_392;

architecture SYN_PLUTO_architecture234 of FD_392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2955 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2955);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture234;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_391 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_391;

architecture SYN_PLUTO_architecture235 of FD_391 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2956 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2956);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture235;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_390 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_390;

architecture SYN_PLUTO_architecture236 of FD_390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2957 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2957);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture236;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_389 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_389;

architecture SYN_PLUTO_architecture237 of FD_389 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2958 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2958);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture237;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_388 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_388;

architecture SYN_PLUTO_architecture238 of FD_388 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2959 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2959);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture238;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_387 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_387;

architecture SYN_PLUTO_architecture239 of FD_387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2960 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2960);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture239;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_386 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_386;

architecture SYN_PLUTO_architecture240 of FD_386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2961 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2961);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture240;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_385 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_385;

architecture SYN_PLUTO_architecture241 of FD_385 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2962 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2962);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture241;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_384 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_384;

architecture SYN_PLUTO_architecture242 of FD_384 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2963 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2963);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture242;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_383 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_383;

architecture SYN_PLUTO_architecture243 of FD_383 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2964 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2964);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture243;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_382 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_382;

architecture SYN_PLUTO_architecture244 of FD_382 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2965 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2965);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture244;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_381 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_381;

architecture SYN_PLUTO_architecture245 of FD_381 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2966 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2966);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture245;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_380 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_380;

architecture SYN_PLUTO_architecture246 of FD_380 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2967 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2967);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture246;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_379 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_379;

architecture SYN_PLUTO_architecture247 of FD_379 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2968 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2968);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture247;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_378 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_378;

architecture SYN_PLUTO_architecture248 of FD_378 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2969 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2969);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture248;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_377 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_377;

architecture SYN_PLUTO of FD_377 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2970 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2970);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_376 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_376;

architecture SYN_PLUTO_architecture of FD_376 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2971 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2971);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_375 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_375;

architecture SYN_PLUTO_architecture2 of FD_375 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2972 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2972);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_374 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_374;

architecture SYN_PLUTO_architecture3 of FD_374 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2973 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2973);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_373 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_373;

architecture SYN_PLUTO_architecture4 of FD_373 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2974 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2974);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_372 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_372;

architecture SYN_PLUTO_architecture5 of FD_372 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2975 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2975);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_371 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_371;

architecture SYN_PLUTO_architecture6 of FD_371 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2976 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2976);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_370 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_370;

architecture SYN_PLUTO_architecture7 of FD_370 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2977 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2977);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_369 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_369;

architecture SYN_PLUTO_architecture8 of FD_369 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2978 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2978);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_368 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_368;

architecture SYN_PLUTO_architecture9 of FD_368 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2979 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2979);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_367 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_367;

architecture SYN_PLUTO_architecture10 of FD_367 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2980 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2980);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_366 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_366;

architecture SYN_PLUTO_architecture11 of FD_366 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2981 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2981);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_365 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_365;

architecture SYN_PLUTO_architecture12 of FD_365 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2982 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2982);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_364 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_364;

architecture SYN_PLUTO_architecture13 of FD_364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2983 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2983);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_363 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_363;

architecture SYN_PLUTO_architecture14 of FD_363 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2984 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2984);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_362 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_362;

architecture SYN_PLUTO_architecture15 of FD_362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2985 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2985);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_361 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_361;

architecture SYN_PLUTO_architecture16 of FD_361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2986 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2986);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_360 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_360;

architecture SYN_PLUTO_architecture17 of FD_360 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2987 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2987);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_359 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_359;

architecture SYN_PLUTO_architecture18 of FD_359 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2988 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2988);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_358 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_358;

architecture SYN_PLUTO_architecture19 of FD_358 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2989 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2989);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_357 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_357;

architecture SYN_PLUTO_architecture20 of FD_357 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2990 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2990);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_356 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_356;

architecture SYN_PLUTO_architecture21 of FD_356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2991 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2991);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_355 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_355;

architecture SYN_PLUTO_architecture22 of FD_355 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2992 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2992);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_354 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_354;

architecture SYN_PLUTO_architecture23 of FD_354 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2993 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2993);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_353 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_353;

architecture SYN_PLUTO_architecture24 of FD_353 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2994 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2994);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_352 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_352;

architecture SYN_PLUTO_architecture25 of FD_352 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2995 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2995);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_351 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_351;

architecture SYN_PLUTO_architecture26 of FD_351 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2996 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2996);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_350 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_350;

architecture SYN_PLUTO_architecture27 of FD_350 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2997 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2997);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_349 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_349;

architecture SYN_PLUTO_architecture28 of FD_349 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2998 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2998);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_348 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_348;

architecture SYN_PLUTO_architecture29 of FD_348 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_2999 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_2999);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_347 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_347;

architecture SYN_PLUTO_architecture30 of FD_347 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3000 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3000);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_346 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_346;

architecture SYN_PLUTO_architecture31 of FD_346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3001 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3001);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_345 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_345;

architecture SYN_PLUTO of FD_345 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3002 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3002);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_344 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_344;

architecture SYN_PLUTO_architecture of FD_344 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3003 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3003);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_343 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_343;

architecture SYN_PLUTO_architecture2 of FD_343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3004 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3004);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_342 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_342;

architecture SYN_PLUTO_architecture3 of FD_342 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3005 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3005);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_341 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_341;

architecture SYN_PLUTO_architecture4 of FD_341 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3006 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3006);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_340 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_340;

architecture SYN_PLUTO_architecture5 of FD_340 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3007 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3007);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_339 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_339;

architecture SYN_PLUTO_architecture6 of FD_339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3008 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3008);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_338 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_338;

architecture SYN_PLUTO_architecture7 of FD_338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3009 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3009);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_337 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_337;

architecture SYN_PLUTO_architecture8 of FD_337 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3010 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3010);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_336 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_336;

architecture SYN_PLUTO_architecture9 of FD_336 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3011 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3011);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_335 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_335;

architecture SYN_PLUTO_architecture10 of FD_335 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3012 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3012);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_334 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_334;

architecture SYN_PLUTO_architecture11 of FD_334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3013 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3013);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_333 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_333;

architecture SYN_PLUTO_architecture12 of FD_333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3014 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3014);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_332 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_332;

architecture SYN_PLUTO_architecture13 of FD_332 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3015 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3015);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_331 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_331;

architecture SYN_PLUTO_architecture14 of FD_331 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3016 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3016);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_330 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_330;

architecture SYN_PLUTO_architecture15 of FD_330 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3017 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3017);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_329 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_329;

architecture SYN_PLUTO_architecture16 of FD_329 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3018 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3018);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_328 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_328;

architecture SYN_PLUTO_architecture17 of FD_328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3019 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3019);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_327 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_327;

architecture SYN_PLUTO_architecture18 of FD_327 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3020 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3020);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_326 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_326;

architecture SYN_PLUTO_architecture19 of FD_326 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3021 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3021);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_325 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_325;

architecture SYN_PLUTO_architecture20 of FD_325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3022 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3022);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_324 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_324;

architecture SYN_PLUTO_architecture21 of FD_324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3023 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3023);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_323 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_323;

architecture SYN_PLUTO_architecture22 of FD_323 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3024 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3024);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_322 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_322;

architecture SYN_PLUTO_architecture23 of FD_322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3025 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3025);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_321 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_321;

architecture SYN_PLUTO_architecture24 of FD_321 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3026 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3026);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_320 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_320;

architecture SYN_PLUTO_architecture25 of FD_320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3027 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3027);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_319 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_319;

architecture SYN_PLUTO_architecture26 of FD_319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3028 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3028);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_318 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_318;

architecture SYN_PLUTO_architecture27 of FD_318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3029 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3029);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_317 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_317;

architecture SYN_PLUTO_architecture28 of FD_317 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3030 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3030);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_316 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_316;

architecture SYN_PLUTO_architecture29 of FD_316 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3031 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3031);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_315 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_315;

architecture SYN_PLUTO_architecture30 of FD_315 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3032 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3032);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_314 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_314;

architecture SYN_PLUTO_architecture31 of FD_314 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3033 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3033);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_313 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_313;

architecture SYN_PLUTO_architecture32 of FD_313 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3034 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3034);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_312 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_312;

architecture SYN_PLUTO_architecture33 of FD_312 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3035 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3035);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_311 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_311;

architecture SYN_PLUTO_architecture34 of FD_311 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3036 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3036);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_310 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_310;

architecture SYN_PLUTO_architecture35 of FD_310 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3037 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3037);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_309 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_309;

architecture SYN_PLUTO_architecture36 of FD_309 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3038 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3038);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_308 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_308;

architecture SYN_PLUTO_architecture37 of FD_308 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3039 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3039);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_307 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_307;

architecture SYN_PLUTO_architecture38 of FD_307 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3040 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3040);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_306 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_306;

architecture SYN_PLUTO_architecture39 of FD_306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3041 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3041);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_305 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_305;

architecture SYN_PLUTO_architecture40 of FD_305 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3042 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3042);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_304 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_304;

architecture SYN_PLUTO_architecture41 of FD_304 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3043 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3043);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_303 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_303;

architecture SYN_PLUTO_architecture42 of FD_303 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3044 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3044);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_302 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_302;

architecture SYN_PLUTO_architecture43 of FD_302 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3045 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3045);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_301 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_301;

architecture SYN_PLUTO_architecture44 of FD_301 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3046 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3046);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_300 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_300;

architecture SYN_PLUTO_architecture45 of FD_300 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3047 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3047);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_299 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_299;

architecture SYN_PLUTO_architecture46 of FD_299 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3048 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3048);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_298 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_298;

architecture SYN_PLUTO_architecture47 of FD_298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3049 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3049);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_297 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_297;

architecture SYN_PLUTO_architecture48 of FD_297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3050 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3050);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_296 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_296;

architecture SYN_PLUTO_architecture49 of FD_296 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3051 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3051);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_295 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_295;

architecture SYN_PLUTO_architecture50 of FD_295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3052 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3052);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_294 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_294;

architecture SYN_PLUTO_architecture51 of FD_294 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3053 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3053);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_293 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_293;

architecture SYN_PLUTO_architecture52 of FD_293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3054 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3054);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_292 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_292;

architecture SYN_PLUTO_architecture53 of FD_292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3055 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3055);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_291 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_291;

architecture SYN_PLUTO_architecture54 of FD_291 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3056 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3056);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_290 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_290;

architecture SYN_PLUTO_architecture55 of FD_290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3057 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3057);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_289 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_289;

architecture SYN_PLUTO_architecture56 of FD_289 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3058 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3058);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_288 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_288;

architecture SYN_PLUTO_architecture57 of FD_288 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3059 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3059);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_287 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_287;

architecture SYN_PLUTO_architecture58 of FD_287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3060 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3060);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_286 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_286;

architecture SYN_PLUTO_architecture59 of FD_286 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3061 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3061);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_285 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_285;

architecture SYN_PLUTO_architecture60 of FD_285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3062 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3062);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_284 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_284;

architecture SYN_PLUTO_architecture61 of FD_284 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3063 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3063);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_283 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_283;

architecture SYN_PLUTO_architecture62 of FD_283 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3064 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3064);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_282 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_282;

architecture SYN_PLUTO_architecture63 of FD_282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3065 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3065);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_281 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_281;

architecture SYN_PLUTO_architecture64 of FD_281 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3066 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3066);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_280 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_280;

architecture SYN_PLUTO_architecture65 of FD_280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3067 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3067);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_279 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_279;

architecture SYN_PLUTO_architecture66 of FD_279 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3068 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3068);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_278 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_278;

architecture SYN_PLUTO_architecture67 of FD_278 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3069 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3069);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_277 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_277;

architecture SYN_PLUTO_architecture68 of FD_277 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3070 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3070);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_276 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_276;

architecture SYN_PLUTO_architecture69 of FD_276 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3071 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3071);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_275 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_275;

architecture SYN_PLUTO_architecture70 of FD_275 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3072 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3072);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_274 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_274;

architecture SYN_PLUTO_architecture71 of FD_274 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3073 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3073);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_273 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_273;

architecture SYN_PLUTO_architecture72 of FD_273 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3074 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3074);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_272 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_272;

architecture SYN_PLUTO_architecture73 of FD_272 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3075 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3075);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_271 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_271;

architecture SYN_PLUTO_architecture74 of FD_271 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3076 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3076);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_270 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_270;

architecture SYN_PLUTO_architecture75 of FD_270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3077 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3077);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_269 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_269;

architecture SYN_PLUTO_architecture76 of FD_269 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3078 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3078);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_268 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_268;

architecture SYN_PLUTO_architecture77 of FD_268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3079 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3079);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_267 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_267;

architecture SYN_PLUTO_architecture78 of FD_267 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3080 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3080);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_266 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_266;

architecture SYN_PLUTO_architecture79 of FD_266 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3081 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3081);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_265 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_265;

architecture SYN_PLUTO_architecture80 of FD_265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3082 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3082);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_264 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_264;

architecture SYN_PLUTO_architecture81 of FD_264 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3083 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3083);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_263 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_263;

architecture SYN_PLUTO_architecture82 of FD_263 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3084 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3084);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_262 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_262;

architecture SYN_PLUTO_architecture83 of FD_262 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3085 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3085);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_261 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_261;

architecture SYN_PLUTO_architecture84 of FD_261 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3086 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3086);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_260 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_260;

architecture SYN_PLUTO_architecture85 of FD_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3087 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3087);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_259 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_259;

architecture SYN_PLUTO_architecture86 of FD_259 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3088 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3088);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_258 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_258;

architecture SYN_PLUTO_architecture87 of FD_258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3089 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3089);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_257 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_257;

architecture SYN_PLUTO_architecture88 of FD_257 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3090 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3090);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_256 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_256;

architecture SYN_PLUTO_architecture89 of FD_256 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3091 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3091);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_255 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_255;

architecture SYN_PLUTO_architecture90 of FD_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3092 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3092);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_254 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_254;

architecture SYN_PLUTO_architecture91 of FD_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3093 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3093);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_253 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_253;

architecture SYN_PLUTO_architecture92 of FD_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3094 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3094);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_252 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_252;

architecture SYN_PLUTO_architecture93 of FD_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3095 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3095);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_251 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_251;

architecture SYN_PLUTO_architecture94 of FD_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3096 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3096);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_250 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_250;

architecture SYN_PLUTO_architecture95 of FD_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3097 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3097);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_249 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_249;

architecture SYN_PLUTO_architecture96 of FD_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3098 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3098);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_248 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_248;

architecture SYN_PLUTO_architecture97 of FD_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3099 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3099);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_247 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_247;

architecture SYN_PLUTO_architecture98 of FD_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3100 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3100);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_246 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_246;

architecture SYN_PLUTO_architecture99 of FD_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3101 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3101);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_245 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_245;

architecture SYN_PLUTO_architecture100 of FD_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3102 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3102);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_244 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_244;

architecture SYN_PLUTO_architecture101 of FD_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3103 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3103);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_243 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_243;

architecture SYN_PLUTO_architecture102 of FD_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3104 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3104);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_242 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_242;

architecture SYN_PLUTO_architecture103 of FD_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3105 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3105);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_241 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_241;

architecture SYN_PLUTO_architecture104 of FD_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3106 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3106);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_240 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_240;

architecture SYN_PLUTO_architecture105 of FD_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3107 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3107);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_239 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_239;

architecture SYN_PLUTO_architecture106 of FD_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3108 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3108);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_238 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_238;

architecture SYN_PLUTO_architecture107 of FD_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3109 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3109);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_237 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_237;

architecture SYN_PLUTO_architecture108 of FD_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3110 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3110);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_236 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_236;

architecture SYN_PLUTO_architecture109 of FD_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3111 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3111);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_235 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_235;

architecture SYN_PLUTO_architecture110 of FD_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3112 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3112);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_234 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_234;

architecture SYN_PLUTO_architecture111 of FD_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3113 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3113);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_233 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_233;

architecture SYN_PLUTO_architecture112 of FD_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3114 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3114);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_232 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_232;

architecture SYN_PLUTO_architecture113 of FD_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3115 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3115);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_231 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_231;

architecture SYN_PLUTO_architecture114 of FD_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3116 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3116);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_230 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_230;

architecture SYN_PLUTO_architecture115 of FD_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3117 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3117);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_229 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_229;

architecture SYN_PLUTO_architecture116 of FD_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3118 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3118);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_228 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_228;

architecture SYN_PLUTO_architecture117 of FD_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3119 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3119);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_227 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_227;

architecture SYN_PLUTO_architecture118 of FD_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3120 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3120);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_226 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_226;

architecture SYN_PLUTO_architecture119 of FD_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3121 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3121);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_225 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_225;

architecture SYN_PLUTO_architecture120 of FD_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3122 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3122);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_224 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_224;

architecture SYN_PLUTO_architecture121 of FD_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3123 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3123);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_223 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_223;

architecture SYN_PLUTO_architecture122 of FD_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3124 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3124);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_222 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_222;

architecture SYN_PLUTO_architecture123 of FD_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3125 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3125);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_221 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_221;

architecture SYN_PLUTO_architecture124 of FD_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3126 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3126);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_220 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_220;

architecture SYN_PLUTO_architecture125 of FD_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3127 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3127);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_219 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_219;

architecture SYN_PLUTO_architecture126 of FD_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3128 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3128);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_218 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_218;

architecture SYN_PLUTO_architecture127 of FD_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3129 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3129);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_217 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_217;

architecture SYN_PLUTO_architecture128 of FD_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3130 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3130);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_216 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_216;

architecture SYN_PLUTO_architecture129 of FD_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3131 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3131);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_215 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_215;

architecture SYN_PLUTO_architecture130 of FD_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3132 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3132);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_214 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_214;

architecture SYN_PLUTO_architecture131 of FD_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3133 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3133);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_213 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_213;

architecture SYN_PLUTO_architecture132 of FD_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3134 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3134);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_212 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_212;

architecture SYN_PLUTO_architecture133 of FD_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3135 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3135);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_211 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_211;

architecture SYN_PLUTO_architecture134 of FD_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3136 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3136);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_210 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_210;

architecture SYN_PLUTO_architecture135 of FD_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3137 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3137);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_209 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_209;

architecture SYN_PLUTO_architecture136 of FD_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3138 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3138);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_208 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_208;

architecture SYN_PLUTO_architecture137 of FD_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3139 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3139);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_207 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_207;

architecture SYN_PLUTO_architecture138 of FD_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3140 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3140);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_206 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_206;

architecture SYN_PLUTO_architecture139 of FD_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3141 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3141);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_205 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_205;

architecture SYN_PLUTO_architecture140 of FD_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3142 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3142);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_204 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_204;

architecture SYN_PLUTO_architecture141 of FD_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3143 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3143);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_203 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_203;

architecture SYN_PLUTO_architecture142 of FD_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3144 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3144);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_202 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_202;

architecture SYN_PLUTO_architecture143 of FD_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3145 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3145);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture143;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_201 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_201;

architecture SYN_PLUTO_architecture144 of FD_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3146 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3146);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture144;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_200 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_200;

architecture SYN_PLUTO_architecture145 of FD_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3147 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3147);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture145;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_199 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_199;

architecture SYN_PLUTO_architecture146 of FD_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3148 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3148);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture146;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_198 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_198;

architecture SYN_PLUTO_architecture147 of FD_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3149 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3149);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture147;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_197 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_197;

architecture SYN_PLUTO_architecture148 of FD_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3150 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3150);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture148;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_196 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_196;

architecture SYN_PLUTO_architecture149 of FD_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3151 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3151);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture149;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_195 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_195;

architecture SYN_PLUTO_architecture150 of FD_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3152 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3152);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture150;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_194 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_194;

architecture SYN_PLUTO_architecture151 of FD_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3153 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3153);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture151;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_193 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_193;

architecture SYN_PLUTO_architecture152 of FD_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3154 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3154);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture152;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_192 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_192;

architecture SYN_PLUTO_architecture153 of FD_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3155 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3155);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture153;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_191 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_191;

architecture SYN_PLUTO_architecture154 of FD_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3156 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3156);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture154;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_190 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_190;

architecture SYN_PLUTO_architecture155 of FD_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3157 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3157);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture155;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_189 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_189;

architecture SYN_PLUTO_architecture156 of FD_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3158 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3158);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture156;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_188 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_188;

architecture SYN_PLUTO_architecture157 of FD_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3159 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3159);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture157;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_187 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_187;

architecture SYN_PLUTO_architecture158 of FD_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3160 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3160);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture158;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_186 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_186;

architecture SYN_PLUTO_architecture159 of FD_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3161 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3161);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture159;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_185 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_185;

architecture SYN_PLUTO_architecture160 of FD_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3162 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3162);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture160;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_184 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_184;

architecture SYN_PLUTO_architecture161 of FD_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3163 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3163);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture161;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_183 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_183;

architecture SYN_PLUTO_architecture162 of FD_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3164 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3164);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture162;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_182 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_182;

architecture SYN_PLUTO_architecture163 of FD_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3165 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3165);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture163;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_181 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_181;

architecture SYN_PLUTO_architecture164 of FD_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3166 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3166);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture164;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_180 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_180;

architecture SYN_PLUTO_architecture165 of FD_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3167 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3167);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture165;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_179 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_179;

architecture SYN_PLUTO_architecture166 of FD_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3168 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3168);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture166;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_178 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_178;

architecture SYN_PLUTO_architecture167 of FD_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3169 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3169);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture167;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_177 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_177;

architecture SYN_PLUTO_architecture168 of FD_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3170 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3170);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture168;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_176 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_176;

architecture SYN_PLUTO_architecture169 of FD_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3171 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3171);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture169;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_175 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_175;

architecture SYN_PLUTO_architecture170 of FD_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3172 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3172);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture170;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_174 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_174;

architecture SYN_PLUTO_architecture171 of FD_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3173 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3173);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture171;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_173 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_173;

architecture SYN_PLUTO_architecture172 of FD_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3174 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3174);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture172;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_172 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_172;

architecture SYN_PLUTO_architecture173 of FD_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3175 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3175);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture173;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_171 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_171;

architecture SYN_PLUTO_architecture174 of FD_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3176 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3176);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture174;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_170 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_170;

architecture SYN_PLUTO_architecture175 of FD_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3177 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3177);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture175;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_169 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_169;

architecture SYN_PLUTO_architecture176 of FD_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3178 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3178);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture176;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_168 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_168;

architecture SYN_PLUTO_architecture177 of FD_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3179 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3179);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture177;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_167 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_167;

architecture SYN_PLUTO_architecture178 of FD_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3180 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3180);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture178;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_166 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_166;

architecture SYN_PLUTO_architecture179 of FD_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3181 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3181);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture179;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_165 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_165;

architecture SYN_PLUTO_architecture180 of FD_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3182 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3182);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture180;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_164 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_164;

architecture SYN_PLUTO_architecture181 of FD_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3183 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3183);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture181;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_163 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_163;

architecture SYN_PLUTO_architecture182 of FD_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3184 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3184);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture182;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_162 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_162;

architecture SYN_PLUTO_architecture183 of FD_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3185 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3185);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture183;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_161 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_161;

architecture SYN_PLUTO_architecture184 of FD_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3186 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3186);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture184;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_160 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_160;

architecture SYN_PLUTO_architecture185 of FD_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3187 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3187);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture185;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_159 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_159;

architecture SYN_PLUTO_architecture186 of FD_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3188 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3188);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture186;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_158 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_158;

architecture SYN_PLUTO_architecture187 of FD_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3189 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3189);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture187;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_157 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_157;

architecture SYN_PLUTO_architecture188 of FD_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3190 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3190);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture188;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_156 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_156;

architecture SYN_PLUTO_architecture189 of FD_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3191 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3191);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture189;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_155 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_155;

architecture SYN_PLUTO_architecture190 of FD_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3192 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3192);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture190;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_154 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_154;

architecture SYN_PLUTO_architecture191 of FD_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3193 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3193);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture191;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_153 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_153;

architecture SYN_PLUTO_architecture192 of FD_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3194 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3194);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture192;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_152 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_152;

architecture SYN_PLUTO_architecture193 of FD_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3195 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3195);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture193;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_151 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_151;

architecture SYN_PLUTO_architecture194 of FD_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3196 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3196);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture194;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_150 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_150;

architecture SYN_PLUTO_architecture195 of FD_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3197 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3197);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture195;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_149 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_149;

architecture SYN_PLUTO_architecture196 of FD_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3198 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3198);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture196;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_148 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_148;

architecture SYN_PLUTO_architecture197 of FD_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3199 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3199);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture197;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_147 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_147;

architecture SYN_PLUTO_architecture198 of FD_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3200 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3200);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture198;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_146 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_146;

architecture SYN_PLUTO_architecture199 of FD_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3201 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3201);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture199;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_145 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_145;

architecture SYN_PLUTO_architecture200 of FD_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3202 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3202);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture200;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_144 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_144;

architecture SYN_PLUTO_architecture201 of FD_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3203 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3203);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture201;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_143 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_143;

architecture SYN_PLUTO_architecture202 of FD_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3204 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3204);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture202;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_142 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_142;

architecture SYN_PLUTO_architecture203 of FD_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3205 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3205);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture203;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_141 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_141;

architecture SYN_PLUTO_architecture204 of FD_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3206 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3206);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture204;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_140 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_140;

architecture SYN_PLUTO_architecture205 of FD_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3207 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3207);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture205;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_139 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_139;

architecture SYN_PLUTO_architecture206 of FD_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3208 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3208);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture206;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_138 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_138;

architecture SYN_PLUTO_architecture207 of FD_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3209 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3209);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture207;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_137 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_137;

architecture SYN_PLUTO_architecture208 of FD_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3210 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3210);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture208;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_136 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_136;

architecture SYN_PLUTO_architecture209 of FD_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3211 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3211);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture209;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_135 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_135;

architecture SYN_PLUTO_architecture210 of FD_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3212 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3212);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture210;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_134 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_134;

architecture SYN_PLUTO_architecture211 of FD_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3213 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3213);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture211;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_133 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_133;

architecture SYN_PLUTO_architecture212 of FD_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3214 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3214);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture212;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_132 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_132;

architecture SYN_PLUTO_architecture213 of FD_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3215 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3215);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture213;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_131 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_131;

architecture SYN_PLUTO_architecture214 of FD_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3216 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3216);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture214;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_130 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_130;

architecture SYN_PLUTO_architecture215 of FD_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3217 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3217);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture215;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_129 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_129;

architecture SYN_PLUTO_architecture216 of FD_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3218 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3218);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture216;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_128 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_128;

architecture SYN_PLUTO_architecture217 of FD_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3219 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3219);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture217;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_127 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_127;

architecture SYN_PLUTO_architecture218 of FD_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3220 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3220);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture218;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_126 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_126;

architecture SYN_PLUTO_architecture219 of FD_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3221 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3221);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture219;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_125 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_125;

architecture SYN_PLUTO_architecture220 of FD_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3222 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3222);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture220;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_124 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_124;

architecture SYN_PLUTO_architecture221 of FD_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3223 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3223);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture221;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_123 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_123;

architecture SYN_PLUTO_architecture222 of FD_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3224 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3224);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture222;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_122 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_122;

architecture SYN_PLUTO_architecture223 of FD_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3225 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3225);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture223;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_121 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_121;

architecture SYN_PLUTO_architecture224 of FD_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3226 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3226);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture224;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_120 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_120;

architecture SYN_PLUTO_architecture225 of FD_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3227 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3227);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture225;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_119 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_119;

architecture SYN_PLUTO_architecture226 of FD_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3228 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3228);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture226;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_118 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_118;

architecture SYN_PLUTO_architecture227 of FD_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3229 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3229);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture227;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_117 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_117;

architecture SYN_PLUTO_architecture228 of FD_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3230 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3230);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture228;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_116 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_116;

architecture SYN_PLUTO_architecture229 of FD_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3231 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3231);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture229;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_115 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_115;

architecture SYN_PLUTO_architecture230 of FD_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3232 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3232);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture230;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_114 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_114;

architecture SYN_PLUTO_architecture231 of FD_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3233 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3233);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture231;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_113 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_113;

architecture SYN_PLUTO_architecture232 of FD_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3234 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3234);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture232;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_112 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_112;

architecture SYN_PLUTO_architecture233 of FD_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3235 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3235);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture233;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_111 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_111;

architecture SYN_PLUTO_architecture234 of FD_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3236 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3236);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture234;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_110 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_110;

architecture SYN_PLUTO_architecture235 of FD_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3237 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3237);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture235;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_109 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_109;

architecture SYN_PLUTO_architecture236 of FD_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3238 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3238);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture236;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_108 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_108;

architecture SYN_PLUTO_architecture237 of FD_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3239 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3239);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture237;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_107 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_107;

architecture SYN_PLUTO_architecture238 of FD_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3240 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3240);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture238;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_106 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_106;

architecture SYN_PLUTO_architecture239 of FD_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3241 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3241);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture239;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_105 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_105;

architecture SYN_PLUTO_architecture240 of FD_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3242 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3242);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture240;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_104 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_104;

architecture SYN_PLUTO_architecture241 of FD_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3243 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3243);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture241;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_103 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_103;

architecture SYN_PLUTO_architecture242 of FD_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3244 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3244);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture242;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_102 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_102;

architecture SYN_PLUTO_architecture243 of FD_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3245 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3245);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture243;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_101 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_101;

architecture SYN_PLUTO_architecture244 of FD_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3246 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3246);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture244;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_100 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_100;

architecture SYN_PLUTO_architecture245 of FD_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3247 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3247);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture245;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_99 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_99;

architecture SYN_PLUTO_architecture246 of FD_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3248 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3248);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture246;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_98 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_98;

architecture SYN_PLUTO_architecture247 of FD_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3249 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3249);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture247;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_97 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_97;

architecture SYN_PLUTO_architecture248 of FD_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3250 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3250);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture248;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_96 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_96;

architecture SYN_PLUTO of FD_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3251 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3251);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_95 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_95;

architecture SYN_PLUTO of FD_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3252 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3252);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_94 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_94;

architecture SYN_PLUTO of FD_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3253 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3253);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_93 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_93;

architecture SYN_PLUTO of FD_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3254 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3254);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_92 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_92;

architecture SYN_PLUTO of FD_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3255 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3255);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_91 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_91;

architecture SYN_PLUTO of FD_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3256 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3256);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_90 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_90;

architecture SYN_PLUTO of FD_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3257 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3257);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_89 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_89;

architecture SYN_PLUTO of FD_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3258 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3258);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_88 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_88;

architecture SYN_PLUTO of FD_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3259 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3259);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_87 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_87;

architecture SYN_PLUTO of FD_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3260 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3260);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_86 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_86;

architecture SYN_PLUTO of FD_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3261 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3261);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_85 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_85;

architecture SYN_PLUTO of FD_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3262 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3262);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_84 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_84;

architecture SYN_PLUTO of FD_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3263 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3263);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_83 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_83;

architecture SYN_PLUTO of FD_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3264 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3264);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_82 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_82;

architecture SYN_PLUTO of FD_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3265 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3265);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_81 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_81;

architecture SYN_PLUTO of FD_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3266 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3266);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_80 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_80;

architecture SYN_PLUTO of FD_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3267 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3267);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_79 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_79;

architecture SYN_PLUTO_architecture of FD_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3268 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3268);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_78 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_78;

architecture SYN_PLUTO_architecture2 of FD_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3269 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3269);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_77 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_77;

architecture SYN_PLUTO_architecture3 of FD_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3270 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3270);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_76 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_76;

architecture SYN_PLUTO_architecture4 of FD_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3271 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3271);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_75 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_75;

architecture SYN_PLUTO_architecture5 of FD_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3272 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3272);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_74 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_74;

architecture SYN_PLUTO_architecture6 of FD_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3273 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3273);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_73 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_73;

architecture SYN_PLUTO_architecture7 of FD_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3274 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3274);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_72 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_72;

architecture SYN_PLUTO_architecture8 of FD_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3275 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3275);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_71 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_71;

architecture SYN_PLUTO_architecture9 of FD_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3276 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3276);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_70 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_70;

architecture SYN_PLUTO_architecture10 of FD_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3277 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3277);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_69 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_69;

architecture SYN_PLUTO_architecture11 of FD_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3278 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3278);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_68 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_68;

architecture SYN_PLUTO_architecture12 of FD_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3279 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3279);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_67 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_67;

architecture SYN_PLUTO_architecture13 of FD_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3280 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3280);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_66 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_66;

architecture SYN_PLUTO_architecture14 of FD_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3281 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3281);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_65 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_65;

architecture SYN_PLUTO_architecture15 of FD_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3282 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3282);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_64 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_64;

architecture SYN_PLUTO of FD_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3283 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3283);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_63 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_63;

architecture SYN_PLUTO_architecture of FD_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3284 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3284);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_62 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_62;

architecture SYN_PLUTO_architecture2 of FD_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3285 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3285);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_61 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_61;

architecture SYN_PLUTO_architecture3 of FD_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3286 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3286);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_60 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_60;

architecture SYN_PLUTO_architecture4 of FD_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3287 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3287);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_59 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_59;

architecture SYN_PLUTO_architecture5 of FD_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3288 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3288);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_58 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_58;

architecture SYN_PLUTO_architecture6 of FD_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3289 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3289);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_57 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_57;

architecture SYN_PLUTO_architecture7 of FD_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3290 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3290);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_56 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_56;

architecture SYN_PLUTO_architecture8 of FD_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3291 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3291);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_55 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_55;

architecture SYN_PLUTO_architecture9 of FD_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3292 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3292);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_54 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_54;

architecture SYN_PLUTO_architecture10 of FD_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3293 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3293);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_53 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_53;

architecture SYN_PLUTO_architecture11 of FD_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3294 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3294);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_52 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_52;

architecture SYN_PLUTO_architecture12 of FD_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3295 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3295);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_51 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_51;

architecture SYN_PLUTO_architecture13 of FD_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3296 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3296);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_50 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_50;

architecture SYN_PLUTO_architecture14 of FD_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3297 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3297);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_49 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_49;

architecture SYN_PLUTO_architecture15 of FD_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3298 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3298);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_48 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_48;

architecture SYN_PLUTO of FD_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3299 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3299);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_47 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_47;

architecture SYN_PLUTO_architecture of FD_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3300 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3300);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_46 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_46;

architecture SYN_PLUTO_architecture2 of FD_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3301 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3301);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_45 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_45;

architecture SYN_PLUTO_architecture3 of FD_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3302 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3302);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_44 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_44;

architecture SYN_PLUTO_architecture4 of FD_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3303 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3303);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_43 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_43;

architecture SYN_PLUTO_architecture5 of FD_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3304 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3304);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_42 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_42;

architecture SYN_PLUTO_architecture6 of FD_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3305 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3305);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_41 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_41;

architecture SYN_PLUTO_architecture7 of FD_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3306 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3306);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_40 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_40;

architecture SYN_PLUTO_architecture8 of FD_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3307 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3307);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_39 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_39;

architecture SYN_PLUTO_architecture9 of FD_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3308 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3308);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_38 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_38;

architecture SYN_PLUTO_architecture10 of FD_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3309 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3309);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_37 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_37;

architecture SYN_PLUTO_architecture11 of FD_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3310 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3310);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_36 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_36;

architecture SYN_PLUTO_architecture12 of FD_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3311 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3311);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_35 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_35;

architecture SYN_PLUTO_architecture13 of FD_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3312 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3312);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_34 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_34;

architecture SYN_PLUTO_architecture14 of FD_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3313 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3313);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_33 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_33;

architecture SYN_PLUTO_architecture15 of FD_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3314 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3314);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_32 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_32;

architecture SYN_PLUTO of FD_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3315 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3315);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_31 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_31;

architecture SYN_PLUTO_architecture of FD_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3316 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3316);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_30 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_30;

architecture SYN_PLUTO_architecture2 of FD_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3317 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3317);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_29 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_29;

architecture SYN_PLUTO_architecture3 of FD_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3318 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3318);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_28 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_28;

architecture SYN_PLUTO_architecture4 of FD_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3319 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3319);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_27 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_27;

architecture SYN_PLUTO_architecture5 of FD_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3320 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3320);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_26 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_26;

architecture SYN_PLUTO_architecture6 of FD_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3321 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3321);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_25 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_25;

architecture SYN_PLUTO_architecture7 of FD_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3322 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3322);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_24 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_24;

architecture SYN_PLUTO_architecture8 of FD_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3323 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3323);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_23 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_23;

architecture SYN_PLUTO_architecture9 of FD_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3324 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3324);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_22 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_22;

architecture SYN_PLUTO_architecture10 of FD_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3325 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3325);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_21 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_21;

architecture SYN_PLUTO_architecture11 of FD_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3326 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3326);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_20 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_20;

architecture SYN_PLUTO_architecture12 of FD_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3327 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3327);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_19 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_19;

architecture SYN_PLUTO_architecture13 of FD_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3328 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3328);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_18 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_18;

architecture SYN_PLUTO_architecture14 of FD_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3329 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3329);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_17 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_17;

architecture SYN_PLUTO_architecture15 of FD_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3330 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3330);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_16 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_16;

architecture SYN_PLUTO of FD_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3331 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3331);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_15 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_15;

architecture SYN_PLUTO_architecture of FD_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3332 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3332);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_14 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_14;

architecture SYN_PLUTO_architecture2 of FD_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3333 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3333);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_13 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_13;

architecture SYN_PLUTO_architecture3 of FD_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3334 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3334);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_12 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_12;

architecture SYN_PLUTO_architecture4 of FD_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3335 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3335);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_11 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_11;

architecture SYN_PLUTO_architecture5 of FD_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3336 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3336);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_10 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_10;

architecture SYN_PLUTO_architecture6 of FD_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3337 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3337);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_9 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_9;

architecture SYN_PLUTO_architecture7 of FD_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3338 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3338);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_8 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_8;

architecture SYN_PLUTO_architecture8 of FD_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3339 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3339);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_7 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_7;

architecture SYN_PLUTO_architecture9 of FD_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3340 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3340);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_6 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_6;

architecture SYN_PLUTO_architecture10 of FD_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3341 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3341);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_5 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_5;

architecture SYN_PLUTO_architecture11 of FD_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3342 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3342);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_4 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_4;

architecture SYN_PLUTO_architecture12 of FD_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3343 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3343);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_3 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_3;

architecture SYN_PLUTO_architecture13 of FD_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3344 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3344);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_2 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_2;

architecture SYN_PLUTO_architecture14 of FD_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3345 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3345);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_1 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_1;

architecture SYN_PLUTO_architecture15 of FD_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_3346 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_3346);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n22_2 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0);  Q 
         : out std_logic_vector (21 downto 0));

end reg_nbit_n22_2;

architecture SYN_struc of reg_nbit_n22_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2207
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2208
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2209
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2210
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2211
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2212
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2213
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2214
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2215
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2216
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2217
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2218
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2219
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2220
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2221
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2222
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2223
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2224
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2225
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2226
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2227
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2228
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   D_I_0 : FD_2228 port map( D => d(0), CK => n2, RESET => reset, Q => Q(0));
   D_I_1 : FD_2227 port map( D => d(1), CK => n2, RESET => reset, Q => Q(1));
   D_I_2 : FD_2226 port map( D => d(2), CK => n2, RESET => reset, Q => Q(2));
   D_I_3 : FD_2225 port map( D => d(3), CK => n2, RESET => reset, Q => Q(3));
   D_I_4 : FD_2224 port map( D => d(4), CK => n2, RESET => reset, Q => Q(4));
   D_I_5 : FD_2223 port map( D => d(5), CK => n2, RESET => reset, Q => Q(5));
   D_I_6 : FD_2222 port map( D => d(6), CK => n2, RESET => reset, Q => Q(6));
   D_I_7 : FD_2221 port map( D => d(7), CK => n2, RESET => reset, Q => Q(7));
   D_I_8 : FD_2220 port map( D => d(8), CK => n2, RESET => reset, Q => Q(8));
   D_I_9 : FD_2219 port map( D => d(9), CK => n2, RESET => reset, Q => Q(9));
   D_I_10 : FD_2218 port map( D => d(10), CK => n2, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2217 port map( D => d(11), CK => n1, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2216 port map( D => d(12), CK => n1, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2215 port map( D => d(13), CK => n1, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2214 port map( D => d(14), CK => n1, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2213 port map( D => d(15), CK => n1, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2212 port map( D => d(16), CK => n1, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2211 port map( D => d(17), CK => n1, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2210 port map( D => d(18), CK => n1, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2209 port map( D => d(19), CK => n1, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2208 port map( D => d(20), CK => n1, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2207 port map( D => d(21), CK => n1, RESET => reset, Q => Q(21))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n2);
   U2 : BUF_X1 port map( A => clk, Z => n1);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n22_1 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0);  Q 
         : out std_logic_vector (21 downto 0));

end reg_nbit_n22_1;

architecture SYN_struc of reg_nbit_n22_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2185
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2186
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2187
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2188
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2189
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2190
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2191
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2192
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2193
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2194
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2195
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2196
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2197
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2198
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2199
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2200
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2201
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2202
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2203
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2204
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2205
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2206
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   D_I_0 : FD_2206 port map( D => d(0), CK => n2, RESET => reset, Q => Q(0));
   D_I_1 : FD_2205 port map( D => d(1), CK => n2, RESET => reset, Q => Q(1));
   D_I_2 : FD_2204 port map( D => d(2), CK => n2, RESET => reset, Q => Q(2));
   D_I_3 : FD_2203 port map( D => d(3), CK => n2, RESET => reset, Q => Q(3));
   D_I_4 : FD_2202 port map( D => d(4), CK => n2, RESET => reset, Q => Q(4));
   D_I_5 : FD_2201 port map( D => d(5), CK => n2, RESET => reset, Q => Q(5));
   D_I_6 : FD_2200 port map( D => d(6), CK => n2, RESET => reset, Q => Q(6));
   D_I_7 : FD_2199 port map( D => d(7), CK => n2, RESET => reset, Q => Q(7));
   D_I_8 : FD_2198 port map( D => d(8), CK => n2, RESET => reset, Q => Q(8));
   D_I_9 : FD_2197 port map( D => d(9), CK => n2, RESET => reset, Q => Q(9));
   D_I_10 : FD_2196 port map( D => d(10), CK => n2, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2195 port map( D => d(11), CK => n1, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2194 port map( D => d(12), CK => n1, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2193 port map( D => d(13), CK => n1, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2192 port map( D => d(14), CK => n1, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2191 port map( D => d(15), CK => n1, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2190 port map( D => d(16), CK => n1, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2189 port map( D => d(17), CK => n1, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2188 port map( D => d(18), CK => n1, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2187 port map( D => d(19), CK => n1, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2186 port map( D => d(20), CK => n1, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2185 port map( D => d(21), CK => n1, RESET => reset, Q => Q(21))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n2);
   U2 : BUF_X1 port map( A => clk, Z => n1);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT8_0 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0);  Co : out std_logic);

end RCA_NBIT8_0;

architecture SYN_STRUCTURAL of RCA_NBIT8_0 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, 
      CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_60 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_59 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_58 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_57 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT8_0 is

   port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (7 downto 0));

end CSB_NBIT8_0;

architecture SYN_STRUCTURAL of CSB_NBIT8_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_NBIT8_7
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT8_0
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_c0_7_port, out_c0_6_port, 
      out_c0_5_port, out_c0_4_port, out_c0_3_port, out_c0_2_port, out_c0_1_port
      , out_c0_0_port, out_c1_7_port, out_c1_6_port, out_c1_5_port, 
      out_c1_4_port, out_c1_3_port, out_c1_2_port, out_c1_1_port, out_c1_0_port
      , n_3347, n_3348 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT8_0 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(7) => 
                           out_c0_7_port, S(6) => out_c0_6_port, S(5) => 
                           out_c0_5_port, S(4) => out_c0_4_port, S(3) => 
                           out_c0_3_port, S(2) => out_c0_2_port, S(1) => 
                           out_c0_1_port, S(0) => out_c0_0_port, Co => n_3347);
   RCA1 : RCA_NBIT8_7 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) 
                           => A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(7) => 
                           out_c1_7_port, S(6) => out_c1_6_port, S(5) => 
                           out_c1_5_port, S(4) => out_c1_4_port, S(3) => 
                           out_c1_3_port, S(2) => out_c1_2_port, S(1) => 
                           out_c1_1_port, S(0) => out_c1_0_port, Co => n_3348);
   U3 : MUX2_X1 port map( A => out_c0_7_port, B => out_c1_7_port, S => Ci, Z =>
                           S(7));
   U4 : MUX2_X1 port map( A => out_c0_6_port, B => out_c1_6_port, S => Ci, Z =>
                           S(6));
   U5 : MUX2_X1 port map( A => out_c0_5_port, B => out_c1_5_port, S => Ci, Z =>
                           S(5));
   U6 : MUX2_X1 port map( A => out_c0_4_port, B => out_c1_4_port, S => Ci, Z =>
                           S(4));
   U7 : MUX2_X1 port map( A => out_c0_3_port, B => out_c1_3_port, S => Ci, Z =>
                           S(3));
   U8 : MUX2_X1 port map( A => out_c0_2_port, B => out_c1_2_port, S => Ci, Z =>
                           S(2));
   U9 : MUX2_X1 port map( A => out_c0_1_port, B => out_c1_1_port, S => Ci, Z =>
                           S(1));
   U10 : MUX2_X1 port map( A => out_c0_0_port, B => out_c1_0_port, S => Ci, Z 
                           => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGSB_0 is

   port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : out
         std_logic);

end PGSB_0;

architecture SYN_BEHAVIORAL of PGSB_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );
   U3 : AND2_X1 port map( A1 => P_in_kj, A2 => P_in_ik, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity GSB_0 is

   port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);

end GSB_0;

architecture SYN_BEHAVIORAL of GSB_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in_ik, B2 => G_in_kj, A => G_in_ik, ZN => n1
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  p, g :
         out std_logic_vector (31 downto 0));

end PG_NBIT32;

architecture SYN_BEHAVIORAL of PG_NBIT32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => p(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => p(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => p(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => p(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => p(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => p(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => p(3));
   U8 : XOR2_X1 port map( A => B(31), B => A(31), Z => p(31));
   U9 : XOR2_X1 port map( A => B(30), B => A(30), Z => p(30));
   U10 : XOR2_X1 port map( A => B(2), B => A(2), Z => p(2));
   U11 : XOR2_X1 port map( A => B(29), B => A(29), Z => p(29));
   U12 : XOR2_X1 port map( A => B(28), B => A(28), Z => p(28));
   U13 : XOR2_X1 port map( A => B(27), B => A(27), Z => p(27));
   U14 : XOR2_X1 port map( A => B(26), B => A(26), Z => p(26));
   U15 : XOR2_X1 port map( A => B(25), B => A(25), Z => p(25));
   U16 : XOR2_X1 port map( A => B(24), B => A(24), Z => p(24));
   U17 : XOR2_X1 port map( A => B(23), B => A(23), Z => p(23));
   U18 : XOR2_X1 port map( A => B(22), B => A(22), Z => p(22));
   U19 : XOR2_X1 port map( A => B(21), B => A(21), Z => p(21));
   U20 : XOR2_X1 port map( A => B(20), B => A(20), Z => p(20));
   U21 : XOR2_X1 port map( A => B(1), B => A(1), Z => p(1));
   U22 : XOR2_X1 port map( A => B(19), B => A(19), Z => p(19));
   U23 : XOR2_X1 port map( A => B(18), B => A(18), Z => p(18));
   U24 : XOR2_X1 port map( A => B(17), B => A(17), Z => p(17));
   U25 : XOR2_X1 port map( A => B(16), B => A(16), Z => p(16));
   U26 : XOR2_X1 port map( A => B(15), B => A(15), Z => p(15));
   U27 : XOR2_X1 port map( A => B(14), B => A(14), Z => p(14));
   U28 : XOR2_X1 port map( A => B(13), B => A(13), Z => p(13));
   U29 : XOR2_X1 port map( A => B(12), B => A(12), Z => p(12));
   U30 : XOR2_X1 port map( A => B(11), B => A(11), Z => p(11));
   U31 : XOR2_X1 port map( A => B(10), B => A(10), Z => p(10));
   U32 : XNOR2_X1 port map( A => n1, B => A(0), ZN => p(0));
   U33 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => g(0));
   U34 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => cin, ZN => n3);
   U35 : INV_X1 port map( A => A(0), ZN => n2);
   U36 : INV_X1 port map( A => B(0), ZN => n1);
   U37 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => g(9));
   U38 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => g(8));
   U39 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => g(7));
   U40 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => g(6));
   U41 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => g(5));
   U42 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => g(4));
   U43 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => g(3));
   U44 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => g(31));
   U45 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => g(30));
   U46 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => g(2));
   U47 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => g(29));
   U48 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => g(28));
   U49 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => g(27));
   U50 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => g(26));
   U51 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => g(25));
   U52 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => g(24));
   U53 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => g(23));
   U54 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => g(22));
   U55 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => g(21));
   U56 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => g(20));
   U57 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => g(1));
   U58 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => g(19));
   U59 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => g(18));
   U60 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => g(17));
   U61 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => g(16));
   U62 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => g(15));
   U63 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => g(14));
   U64 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => g(13));
   U65 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => g(12));
   U66 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => g(11));
   U67 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => g(10));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n16_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0);  Q 
         : out std_logic_vector (15 downto 0));

end reg_nbit_n16_0;

architecture SYN_struc of reg_nbit_n16_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_81
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_82
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_83
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_84
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_85
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_86
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_87
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_88
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_89
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_90
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_91
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_92
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_93
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_94
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_95
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_96
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   D_I_0 : FD_96 port map( D => d(0), CK => n4, RESET => n2, Q => Q(0));
   D_I_1 : FD_95 port map( D => d(1), CK => n4, RESET => n2, Q => Q(1));
   D_I_2 : FD_94 port map( D => d(2), CK => n4, RESET => n2, Q => Q(2));
   D_I_3 : FD_93 port map( D => d(3), CK => n4, RESET => n2, Q => Q(3));
   D_I_4 : FD_92 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_91 port map( D => d(5), CK => n3, RESET => n1, Q => Q(5));
   D_I_6 : FD_90 port map( D => d(6), CK => n3, RESET => n1, Q => Q(6));
   D_I_7 : FD_89 port map( D => d(7), CK => n3, RESET => n1, Q => Q(7));
   D_I_8 : FD_88 port map( D => d(8), CK => n3, RESET => n1, Q => Q(8));
   D_I_9 : FD_87 port map( D => d(9), CK => n3, RESET => n1, Q => Q(9));
   D_I_10 : FD_86 port map( D => d(10), CK => n3, RESET => n1, Q => Q(10));
   D_I_11 : FD_85 port map( D => d(11), CK => n3, RESET => n1, Q => Q(11));
   D_I_12 : FD_84 port map( D => d(12), CK => n3, RESET => n1, Q => Q(12));
   D_I_13 : FD_83 port map( D => d(13), CK => n3, RESET => n1, Q => Q(13));
   D_I_14 : FD_82 port map( D => d(14), CK => n3, RESET => n1, Q => Q(14));
   D_I_15 : FD_81 port map( D => d(15), CK => n3, RESET => n1, Q => Q(15));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT31 is

   port( a, b : in std_logic_vector (30 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (31 downto 0));

end adder_NBIT31;

architecture SYN_beh of adder_NBIT31 is

   component adder_NBIT31_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3349 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT31_DW01_add_0 port map( A(31) => a(30), 
                           A(30) => a(30), A(29) => a(29), A(28) => a(28), 
                           A(27) => a(27), A(26) => a(26), A(25) => a(25), 
                           A(24) => a(24), A(23) => a(23), A(22) => a(22), 
                           A(21) => a(21), A(20) => a(20), A(19) => a(19), 
                           A(18) => a(18), A(17) => a(17), A(16) => a(16), 
                           A(15) => a(15), A(14) => a(14), A(13) => a(13), 
                           A(12) => a(12), A(11) => a(11), A(10) => a(10), A(9)
                           => a(9), A(8) => a(8), A(7) => a(7), A(6) => a(6), 
                           A(5) => a(5), A(4) => a(4), A(3) => a(3), A(2) => 
                           a(2), A(1) => a(1), A(0) => a(0), B(31) => b(30), 
                           B(30) => b(30), B(29) => b(29), B(28) => b(28), 
                           B(27) => b(27), B(26) => b(26), B(25) => b(25), 
                           B(24) => b(24), B(23) => b(23), B(22) => b(22), 
                           B(21) => b(21), B(20) => b(20), B(19) => b(19), 
                           B(18) => b(18), B(17) => b(17), B(16) => b(16), 
                           B(15) => b(15), B(14) => b(14), B(13) => b(13), 
                           B(12) => b(12), B(11) => b(11), B(10) => b(10), B(9)
                           => b(9), B(8) => b(8), B(7) => b(7), B(6) => b(6), 
                           B(5) => b(5), B(4) => b(4), B(3) => b(3), B(2) => 
                           b(2), B(1) => b(1), B(0) => b(0), CI => cin, SUM(31)
                           => s(31), SUM(30) => s(30), SUM(29) => s(29), 
                           SUM(28) => s(28), SUM(27) => s(27), SUM(26) => s(26)
                           , SUM(25) => s(25), SUM(24) => s(24), SUM(23) => 
                           s(23), SUM(22) => s(22), SUM(21) => s(21), SUM(20) 
                           => s(20), SUM(19) => s(19), SUM(18) => s(18), 
                           SUM(17) => s(17), SUM(16) => s(16), SUM(15) => s(15)
                           , SUM(14) => s(14), SUM(13) => s(13), SUM(12) => 
                           s(12), SUM(11) => s(11), SUM(10) => s(10), SUM(9) =>
                           s(9), SUM(8) => s(8), SUM(7) => s(7), SUM(6) => s(6)
                           , SUM(5) => s(5), SUM(4) => s(4), SUM(3) => s(3), 
                           SUM(2) => s(2), SUM(1) => s(1), SUM(0) => s(0), CO 
                           => n_3349);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N31_Z3 is

   port( inputs : in std_logic_vector (0 to 247);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (30 downto 0));

end MUX_zbit_nbit_N31_Z3;

architecture SYN_beh of MUX_zbit_nbit_N31_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, 
      N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, 
      N230, N231, N232, N233, N234, N235, N236, N237, n4, n1, n2, n3, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145 : std_logic;

begin
   
   Y_reg_30_inst : DLH_X1 port map( G => n4, D => N237, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n4, D => N236, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n4, D => N235, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n4, D => N234, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n4, D => N233, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n4, D => N232, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n4, D => N231, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n4, D => N230, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n4, D => N229, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n4, D => N228, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N227, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N226, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N225, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N224, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N223, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N222, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N221, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N220, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N219, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N218, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N217, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N216, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N215, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N214, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N213, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N212, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N211, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N210, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N209, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N208, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N207, Q => Y(0));
   n4 <= '1';
   U3 : OR4_X1 port map( A1 => n10, A2 => n5, A3 => n9, A4 => n142, ZN => n1);
   U4 : INV_X2 port map( A => n1, ZN => n2);
   U5 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n143, ZN => n21);
   U6 : INV_X2 port map( A => n21, ZN => n3);
   U7 : OR3_X1 port map( A1 => n145, A2 => SEL(2), A3 => n144, ZN => n17);
   U8 : INV_X2 port map( A => n17, ZN => n5);
   U9 : OR3_X1 port map( A1 => n143, A2 => SEL(1), A3 => n145, ZN => n19);
   U10 : INV_X2 port map( A => n19, ZN => n6);
   U11 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n144, ZN => n18);
   U12 : INV_X2 port map( A => n18, ZN => n7);
   U13 : OR3_X1 port map( A1 => n145, A2 => n143, A3 => n144, ZN => n20);
   U14 : INV_X2 port map( A => n20, ZN => n8);
   U15 : OR3_X1 port map( A1 => n143, A2 => SEL(0), A3 => n144, ZN => n15);
   U16 : INV_X2 port map( A => n15, ZN => n9);
   U17 : OR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n145, ZN => n16);
   U18 : INV_X2 port map( A => n16, ZN => n10);
   U19 : NAND4_X1 port map( A1 => n11, A2 => n12, A3 => n13, A4 => n14, ZN => 
                           N237);
   U20 : AOI22_X1 port map( A1 => inputs(0), A2 => n2, B1 => inputs(186), B2 =>
                           n9, ZN => n14);
   U21 : AOI22_X1 port map( A1 => inputs(31), A2 => n10, B1 => inputs(93), B2 
                           => n5, ZN => n13);
   U22 : AOI22_X1 port map( A1 => inputs(62), A2 => n7, B1 => inputs(155), B2 
                           => n6, ZN => n12);
   U23 : AOI22_X1 port map( A1 => inputs(217), A2 => n8, B1 => inputs(124), B2 
                           => n3, ZN => n11);
   U24 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           N236);
   U25 : AOI22_X1 port map( A1 => inputs(1), A2 => n2, B1 => inputs(187), B2 =>
                           n9, ZN => n25);
   U26 : AOI22_X1 port map( A1 => inputs(32), A2 => n10, B1 => inputs(94), B2 
                           => n5, ZN => n24);
   U27 : AOI22_X1 port map( A1 => inputs(63), A2 => n7, B1 => inputs(156), B2 
                           => n6, ZN => n23);
   U28 : AOI22_X1 port map( A1 => inputs(218), A2 => n8, B1 => inputs(125), B2 
                           => n3, ZN => n22);
   U29 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n28, A4 => n29, ZN => 
                           N235);
   U30 : AOI22_X1 port map( A1 => inputs(2), A2 => n2, B1 => inputs(188), B2 =>
                           n9, ZN => n29);
   U31 : AOI22_X1 port map( A1 => inputs(33), A2 => n10, B1 => inputs(95), B2 
                           => n5, ZN => n28);
   U32 : AOI22_X1 port map( A1 => inputs(64), A2 => n7, B1 => inputs(157), B2 
                           => n6, ZN => n27);
   U33 : AOI22_X1 port map( A1 => inputs(219), A2 => n8, B1 => inputs(126), B2 
                           => n3, ZN => n26);
   U34 : NAND4_X1 port map( A1 => n30, A2 => n31, A3 => n32, A4 => n33, ZN => 
                           N234);
   U35 : AOI22_X1 port map( A1 => inputs(3), A2 => n2, B1 => inputs(189), B2 =>
                           n9, ZN => n33);
   U36 : AOI22_X1 port map( A1 => inputs(34), A2 => n10, B1 => inputs(96), B2 
                           => n5, ZN => n32);
   U37 : AOI22_X1 port map( A1 => inputs(65), A2 => n7, B1 => inputs(158), B2 
                           => n6, ZN => n31);
   U38 : AOI22_X1 port map( A1 => inputs(220), A2 => n8, B1 => inputs(127), B2 
                           => n3, ZN => n30);
   U39 : NAND4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           N233);
   U40 : AOI22_X1 port map( A1 => inputs(4), A2 => n2, B1 => inputs(190), B2 =>
                           n9, ZN => n37);
   U41 : AOI22_X1 port map( A1 => inputs(35), A2 => n10, B1 => inputs(97), B2 
                           => n5, ZN => n36);
   U42 : AOI22_X1 port map( A1 => inputs(66), A2 => n7, B1 => inputs(159), B2 
                           => n6, ZN => n35);
   U43 : AOI22_X1 port map( A1 => inputs(221), A2 => n8, B1 => inputs(128), B2 
                           => n3, ZN => n34);
   U44 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           N232);
   U45 : AOI22_X1 port map( A1 => inputs(5), A2 => n2, B1 => inputs(191), B2 =>
                           n9, ZN => n41);
   U46 : AOI22_X1 port map( A1 => inputs(36), A2 => n10, B1 => inputs(98), B2 
                           => n5, ZN => n40);
   U47 : AOI22_X1 port map( A1 => inputs(67), A2 => n7, B1 => inputs(160), B2 
                           => n6, ZN => n39);
   U48 : AOI22_X1 port map( A1 => inputs(222), A2 => n8, B1 => inputs(129), B2 
                           => n3, ZN => n38);
   U49 : NAND4_X1 port map( A1 => n42, A2 => n43, A3 => n44, A4 => n45, ZN => 
                           N231);
   U50 : AOI22_X1 port map( A1 => inputs(6), A2 => n2, B1 => inputs(192), B2 =>
                           n9, ZN => n45);
   U51 : AOI22_X1 port map( A1 => inputs(37), A2 => n10, B1 => inputs(99), B2 
                           => n5, ZN => n44);
   U52 : AOI22_X1 port map( A1 => inputs(68), A2 => n7, B1 => inputs(161), B2 
                           => n6, ZN => n43);
   U53 : AOI22_X1 port map( A1 => inputs(223), A2 => n8, B1 => inputs(130), B2 
                           => n3, ZN => n42);
   U54 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           N230);
   U55 : AOI22_X1 port map( A1 => inputs(7), A2 => n2, B1 => inputs(193), B2 =>
                           n9, ZN => n49);
   U56 : AOI22_X1 port map( A1 => inputs(38), A2 => n10, B1 => inputs(100), B2 
                           => n5, ZN => n48);
   U57 : AOI22_X1 port map( A1 => inputs(69), A2 => n7, B1 => inputs(162), B2 
                           => n6, ZN => n47);
   U58 : AOI22_X1 port map( A1 => inputs(224), A2 => n8, B1 => inputs(131), B2 
                           => n3, ZN => n46);
   U59 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           N229);
   U60 : AOI22_X1 port map( A1 => inputs(8), A2 => n2, B1 => inputs(194), B2 =>
                           n9, ZN => n53);
   U61 : AOI22_X1 port map( A1 => inputs(39), A2 => n10, B1 => inputs(101), B2 
                           => n5, ZN => n52);
   U62 : AOI22_X1 port map( A1 => inputs(70), A2 => n7, B1 => inputs(163), B2 
                           => n6, ZN => n51);
   U63 : AOI22_X1 port map( A1 => inputs(225), A2 => n8, B1 => inputs(132), B2 
                           => n3, ZN => n50);
   U64 : NAND4_X1 port map( A1 => n54, A2 => n55, A3 => n56, A4 => n57, ZN => 
                           N228);
   U65 : AOI22_X1 port map( A1 => inputs(9), A2 => n2, B1 => inputs(195), B2 =>
                           n9, ZN => n57);
   U66 : AOI22_X1 port map( A1 => inputs(40), A2 => n10, B1 => inputs(102), B2 
                           => n5, ZN => n56);
   U67 : AOI22_X1 port map( A1 => inputs(71), A2 => n7, B1 => inputs(164), B2 
                           => n6, ZN => n55);
   U68 : AOI22_X1 port map( A1 => inputs(226), A2 => n8, B1 => inputs(133), B2 
                           => n3, ZN => n54);
   U69 : NAND4_X1 port map( A1 => n58, A2 => n59, A3 => n60, A4 => n61, ZN => 
                           N227);
   U70 : AOI22_X1 port map( A1 => inputs(10), A2 => n2, B1 => inputs(196), B2 
                           => n9, ZN => n61);
   U71 : AOI22_X1 port map( A1 => inputs(41), A2 => n10, B1 => inputs(103), B2 
                           => n5, ZN => n60);
   U72 : AOI22_X1 port map( A1 => inputs(72), A2 => n7, B1 => inputs(165), B2 
                           => n6, ZN => n59);
   U73 : AOI22_X1 port map( A1 => inputs(227), A2 => n8, B1 => inputs(134), B2 
                           => n3, ZN => n58);
   U74 : NAND4_X1 port map( A1 => n62, A2 => n63, A3 => n64, A4 => n65, ZN => 
                           N226);
   U75 : AOI22_X1 port map( A1 => inputs(11), A2 => n2, B1 => inputs(197), B2 
                           => n9, ZN => n65);
   U76 : AOI22_X1 port map( A1 => inputs(42), A2 => n10, B1 => inputs(104), B2 
                           => n5, ZN => n64);
   U77 : AOI22_X1 port map( A1 => inputs(73), A2 => n7, B1 => inputs(166), B2 
                           => n6, ZN => n63);
   U78 : AOI22_X1 port map( A1 => inputs(228), A2 => n8, B1 => inputs(135), B2 
                           => n3, ZN => n62);
   U79 : NAND4_X1 port map( A1 => n66, A2 => n67, A3 => n68, A4 => n69, ZN => 
                           N225);
   U80 : AOI22_X1 port map( A1 => inputs(12), A2 => n2, B1 => inputs(198), B2 
                           => n9, ZN => n69);
   U81 : AOI22_X1 port map( A1 => inputs(43), A2 => n10, B1 => inputs(105), B2 
                           => n5, ZN => n68);
   U82 : AOI22_X1 port map( A1 => inputs(74), A2 => n7, B1 => inputs(167), B2 
                           => n6, ZN => n67);
   U83 : AOI22_X1 port map( A1 => inputs(229), A2 => n8, B1 => inputs(136), B2 
                           => n3, ZN => n66);
   U84 : NAND4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           N224);
   U85 : AOI22_X1 port map( A1 => inputs(13), A2 => n2, B1 => inputs(199), B2 
                           => n9, ZN => n73);
   U86 : AOI22_X1 port map( A1 => inputs(44), A2 => n10, B1 => inputs(106), B2 
                           => n5, ZN => n72);
   U87 : AOI22_X1 port map( A1 => inputs(75), A2 => n7, B1 => inputs(168), B2 
                           => n6, ZN => n71);
   U88 : AOI22_X1 port map( A1 => inputs(230), A2 => n8, B1 => inputs(137), B2 
                           => n3, ZN => n70);
   U89 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           N223);
   U90 : AOI22_X1 port map( A1 => inputs(14), A2 => n2, B1 => inputs(200), B2 
                           => n9, ZN => n77);
   U91 : AOI22_X1 port map( A1 => inputs(45), A2 => n10, B1 => inputs(107), B2 
                           => n5, ZN => n76);
   U92 : AOI22_X1 port map( A1 => inputs(76), A2 => n7, B1 => inputs(169), B2 
                           => n6, ZN => n75);
   U93 : AOI22_X1 port map( A1 => inputs(231), A2 => n8, B1 => inputs(138), B2 
                           => n3, ZN => n74);
   U94 : NAND4_X1 port map( A1 => n78, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           N222);
   U95 : AOI22_X1 port map( A1 => inputs(15), A2 => n2, B1 => inputs(201), B2 
                           => n9, ZN => n81);
   U96 : AOI22_X1 port map( A1 => inputs(46), A2 => n10, B1 => inputs(108), B2 
                           => n5, ZN => n80);
   U97 : AOI22_X1 port map( A1 => inputs(77), A2 => n7, B1 => inputs(170), B2 
                           => n6, ZN => n79);
   U98 : AOI22_X1 port map( A1 => inputs(232), A2 => n8, B1 => inputs(139), B2 
                           => n3, ZN => n78);
   U99 : NAND4_X1 port map( A1 => n82, A2 => n83, A3 => n84, A4 => n85, ZN => 
                           N221);
   U100 : AOI22_X1 port map( A1 => inputs(16), A2 => n2, B1 => inputs(202), B2 
                           => n9, ZN => n85);
   U101 : AOI22_X1 port map( A1 => inputs(47), A2 => n10, B1 => inputs(109), B2
                           => n5, ZN => n84);
   U102 : AOI22_X1 port map( A1 => inputs(78), A2 => n7, B1 => inputs(171), B2 
                           => n6, ZN => n83);
   U103 : AOI22_X1 port map( A1 => inputs(233), A2 => n8, B1 => inputs(140), B2
                           => n3, ZN => n82);
   U104 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           N220);
   U105 : AOI22_X1 port map( A1 => inputs(17), A2 => n2, B1 => inputs(203), B2 
                           => n9, ZN => n89);
   U106 : AOI22_X1 port map( A1 => inputs(48), A2 => n10, B1 => inputs(110), B2
                           => n5, ZN => n88);
   U107 : AOI22_X1 port map( A1 => inputs(79), A2 => n7, B1 => inputs(172), B2 
                           => n6, ZN => n87);
   U108 : AOI22_X1 port map( A1 => inputs(234), A2 => n8, B1 => inputs(141), B2
                           => n3, ZN => n86);
   U109 : NAND4_X1 port map( A1 => n90, A2 => n91, A3 => n92, A4 => n93, ZN => 
                           N219);
   U110 : AOI22_X1 port map( A1 => inputs(18), A2 => n2, B1 => inputs(204), B2 
                           => n9, ZN => n93);
   U111 : AOI22_X1 port map( A1 => inputs(49), A2 => n10, B1 => inputs(111), B2
                           => n5, ZN => n92);
   U112 : AOI22_X1 port map( A1 => inputs(80), A2 => n7, B1 => inputs(173), B2 
                           => n6, ZN => n91);
   U113 : AOI22_X1 port map( A1 => inputs(235), A2 => n8, B1 => inputs(142), B2
                           => n3, ZN => n90);
   U114 : NAND4_X1 port map( A1 => n94, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           N218);
   U115 : AOI22_X1 port map( A1 => inputs(19), A2 => n2, B1 => inputs(205), B2 
                           => n9, ZN => n97);
   U116 : AOI22_X1 port map( A1 => inputs(50), A2 => n10, B1 => inputs(112), B2
                           => n5, ZN => n96);
   U117 : AOI22_X1 port map( A1 => inputs(81), A2 => n7, B1 => inputs(174), B2 
                           => n6, ZN => n95);
   U118 : AOI22_X1 port map( A1 => inputs(236), A2 => n8, B1 => inputs(143), B2
                           => n3, ZN => n94);
   U119 : NAND4_X1 port map( A1 => n98, A2 => n99, A3 => n100, A4 => n101, ZN 
                           => N217);
   U120 : AOI22_X1 port map( A1 => inputs(20), A2 => n2, B1 => inputs(206), B2 
                           => n9, ZN => n101);
   U121 : AOI22_X1 port map( A1 => inputs(51), A2 => n10, B1 => inputs(113), B2
                           => n5, ZN => n100);
   U122 : AOI22_X1 port map( A1 => inputs(82), A2 => n7, B1 => inputs(175), B2 
                           => n6, ZN => n99);
   U123 : AOI22_X1 port map( A1 => inputs(237), A2 => n8, B1 => inputs(144), B2
                           => n3, ZN => n98);
   U124 : NAND4_X1 port map( A1 => n102, A2 => n103, A3 => n104, A4 => n105, ZN
                           => N216);
   U125 : AOI22_X1 port map( A1 => inputs(21), A2 => n2, B1 => inputs(207), B2 
                           => n9, ZN => n105);
   U126 : AOI22_X1 port map( A1 => inputs(52), A2 => n10, B1 => inputs(114), B2
                           => n5, ZN => n104);
   U127 : AOI22_X1 port map( A1 => inputs(83), A2 => n7, B1 => inputs(176), B2 
                           => n6, ZN => n103);
   U128 : AOI22_X1 port map( A1 => inputs(238), A2 => n8, B1 => inputs(145), B2
                           => n3, ZN => n102);
   U129 : NAND4_X1 port map( A1 => n106, A2 => n107, A3 => n108, A4 => n109, ZN
                           => N215);
   U130 : AOI22_X1 port map( A1 => inputs(22), A2 => n2, B1 => inputs(208), B2 
                           => n9, ZN => n109);
   U131 : AOI22_X1 port map( A1 => inputs(53), A2 => n10, B1 => inputs(115), B2
                           => n5, ZN => n108);
   U132 : AOI22_X1 port map( A1 => inputs(84), A2 => n7, B1 => inputs(177), B2 
                           => n6, ZN => n107);
   U133 : AOI22_X1 port map( A1 => inputs(239), A2 => n8, B1 => inputs(146), B2
                           => n3, ZN => n106);
   U134 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN
                           => N214);
   U135 : AOI22_X1 port map( A1 => inputs(23), A2 => n2, B1 => inputs(209), B2 
                           => n9, ZN => n113);
   U136 : AOI22_X1 port map( A1 => inputs(54), A2 => n10, B1 => inputs(116), B2
                           => n5, ZN => n112);
   U137 : AOI22_X1 port map( A1 => inputs(85), A2 => n7, B1 => inputs(178), B2 
                           => n6, ZN => n111);
   U138 : AOI22_X1 port map( A1 => inputs(240), A2 => n8, B1 => inputs(147), B2
                           => n3, ZN => n110);
   U139 : NAND4_X1 port map( A1 => n114, A2 => n115, A3 => n116, A4 => n117, ZN
                           => N213);
   U140 : AOI22_X1 port map( A1 => inputs(24), A2 => n2, B1 => inputs(210), B2 
                           => n9, ZN => n117);
   U141 : AOI22_X1 port map( A1 => inputs(55), A2 => n10, B1 => inputs(117), B2
                           => n5, ZN => n116);
   U142 : AOI22_X1 port map( A1 => inputs(86), A2 => n7, B1 => inputs(179), B2 
                           => n6, ZN => n115);
   U143 : AOI22_X1 port map( A1 => inputs(241), A2 => n8, B1 => inputs(148), B2
                           => n3, ZN => n114);
   U144 : NAND4_X1 port map( A1 => n118, A2 => n119, A3 => n120, A4 => n121, ZN
                           => N212);
   U145 : AOI22_X1 port map( A1 => inputs(25), A2 => n2, B1 => inputs(211), B2 
                           => n9, ZN => n121);
   U146 : AOI22_X1 port map( A1 => inputs(56), A2 => n10, B1 => inputs(118), B2
                           => n5, ZN => n120);
   U147 : AOI22_X1 port map( A1 => inputs(87), A2 => n7, B1 => inputs(180), B2 
                           => n6, ZN => n119);
   U148 : AOI22_X1 port map( A1 => inputs(242), A2 => n8, B1 => inputs(149), B2
                           => n3, ZN => n118);
   U149 : NAND4_X1 port map( A1 => n122, A2 => n123, A3 => n124, A4 => n125, ZN
                           => N211);
   U150 : AOI22_X1 port map( A1 => inputs(26), A2 => n2, B1 => inputs(212), B2 
                           => n9, ZN => n125);
   U151 : AOI22_X1 port map( A1 => inputs(57), A2 => n10, B1 => inputs(119), B2
                           => n5, ZN => n124);
   U152 : AOI22_X1 port map( A1 => inputs(88), A2 => n7, B1 => inputs(181), B2 
                           => n6, ZN => n123);
   U153 : AOI22_X1 port map( A1 => inputs(243), A2 => n8, B1 => inputs(150), B2
                           => n3, ZN => n122);
   U154 : NAND4_X1 port map( A1 => n126, A2 => n127, A3 => n128, A4 => n129, ZN
                           => N210);
   U155 : AOI22_X1 port map( A1 => inputs(27), A2 => n2, B1 => inputs(213), B2 
                           => n9, ZN => n129);
   U156 : AOI22_X1 port map( A1 => inputs(58), A2 => n10, B1 => inputs(120), B2
                           => n5, ZN => n128);
   U157 : AOI22_X1 port map( A1 => inputs(89), A2 => n7, B1 => inputs(182), B2 
                           => n6, ZN => n127);
   U158 : AOI22_X1 port map( A1 => inputs(244), A2 => n8, B1 => inputs(151), B2
                           => n3, ZN => n126);
   U159 : NAND4_X1 port map( A1 => n130, A2 => n131, A3 => n132, A4 => n133, ZN
                           => N209);
   U160 : AOI22_X1 port map( A1 => inputs(28), A2 => n2, B1 => inputs(214), B2 
                           => n9, ZN => n133);
   U161 : AOI22_X1 port map( A1 => inputs(59), A2 => n10, B1 => inputs(121), B2
                           => n5, ZN => n132);
   U162 : AOI22_X1 port map( A1 => inputs(90), A2 => n7, B1 => inputs(183), B2 
                           => n6, ZN => n131);
   U163 : AOI22_X1 port map( A1 => inputs(245), A2 => n8, B1 => inputs(152), B2
                           => n3, ZN => n130);
   U164 : NAND4_X1 port map( A1 => n134, A2 => n135, A3 => n136, A4 => n137, ZN
                           => N208);
   U165 : AOI22_X1 port map( A1 => inputs(29), A2 => n2, B1 => inputs(215), B2 
                           => n9, ZN => n137);
   U166 : AOI22_X1 port map( A1 => inputs(60), A2 => n10, B1 => inputs(122), B2
                           => n5, ZN => n136);
   U167 : AOI22_X1 port map( A1 => inputs(91), A2 => n7, B1 => inputs(184), B2 
                           => n6, ZN => n135);
   U168 : AOI22_X1 port map( A1 => inputs(246), A2 => n8, B1 => inputs(153), B2
                           => n3, ZN => n134);
   U169 : NAND4_X1 port map( A1 => n138, A2 => n139, A3 => n140, A4 => n141, ZN
                           => N207);
   U171 : AOI22_X1 port map( A1 => inputs(30), A2 => n2, B1 => inputs(216), B2 
                           => n9, ZN => n141);
   U172 : OR4_X1 port map( A1 => n3, A2 => n8, A3 => n6, A4 => n7, ZN => n142);
   U173 : AOI22_X1 port map( A1 => inputs(61), A2 => n10, B1 => inputs(123), B2
                           => n5, ZN => n140);
   U174 : AOI22_X1 port map( A1 => inputs(92), A2 => n7, B1 => inputs(185), B2 
                           => n6, ZN => n139);
   U175 : AOI22_X1 port map( A1 => inputs(247), A2 => n8, B1 => inputs(154), B2
                           => n3, ZN => n138);
   U176 : INV_X1 port map( A => SEL(1), ZN => n144);
   U177 : INV_X1 port map( A => SEL(2), ZN => n143);
   U178 : INV_X1 port map( A => SEL(0), ZN => n145);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT29 is

   port( a, b : in std_logic_vector (28 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (29 downto 0));

end adder_NBIT29;

architecture SYN_beh of adder_NBIT29 is

   component adder_NBIT29_DW01_add_0
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3350 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT29_DW01_add_0 port map( A(29) => a(28), 
                           A(28) => a(28), A(27) => a(27), A(26) => a(26), 
                           A(25) => a(25), A(24) => a(24), A(23) => a(23), 
                           A(22) => a(22), A(21) => a(21), A(20) => a(20), 
                           A(19) => a(19), A(18) => a(18), A(17) => a(17), 
                           A(16) => a(16), A(15) => a(15), A(14) => a(14), 
                           A(13) => a(13), A(12) => a(12), A(11) => a(11), 
                           A(10) => a(10), A(9) => a(9), A(8) => a(8), A(7) => 
                           a(7), A(6) => a(6), A(5) => a(5), A(4) => a(4), A(3)
                           => a(3), A(2) => a(2), A(1) => a(1), A(0) => a(0), 
                           B(29) => b(28), B(28) => b(28), B(27) => b(27), 
                           B(26) => b(26), B(25) => b(25), B(24) => b(24), 
                           B(23) => b(23), B(22) => b(22), B(21) => b(21), 
                           B(20) => b(20), B(19) => b(19), B(18) => b(18), 
                           B(17) => b(17), B(16) => b(16), B(15) => b(15), 
                           B(14) => b(14), B(13) => b(13), B(12) => b(12), 
                           B(11) => b(11), B(10) => b(10), B(9) => b(9), B(8) 
                           => b(8), B(7) => b(7), B(6) => b(6), B(5) => b(5), 
                           B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1) => 
                           b(1), B(0) => b(0), CI => cin, SUM(29) => s(29), 
                           SUM(28) => s(28), SUM(27) => s(27), SUM(26) => s(26)
                           , SUM(25) => s(25), SUM(24) => s(24), SUM(23) => 
                           s(23), SUM(22) => s(22), SUM(21) => s(21), SUM(20) 
                           => s(20), SUM(19) => s(19), SUM(18) => s(18), 
                           SUM(17) => s(17), SUM(16) => s(16), SUM(15) => s(15)
                           , SUM(14) => s(14), SUM(13) => s(13), SUM(12) => 
                           s(12), SUM(11) => s(11), SUM(10) => s(10), SUM(9) =>
                           s(9), SUM(8) => s(8), SUM(7) => s(7), SUM(6) => s(6)
                           , SUM(5) => s(5), SUM(4) => s(4), SUM(3) => s(3), 
                           SUM(2) => s(2), SUM(1) => s(1), SUM(0) => s(0), CO 
                           => n_3350);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N29_Z3 is

   port( inputs : in std_logic_vector (0 to 231);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (28 downto 0));

end MUX_zbit_nbit_N29_Z3;

architecture SYN_beh of MUX_zbit_nbit_N29_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, 
      N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, 
      N218, N219, N220, N221, N222, N223, n4, n1, n2, n3, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137 : std_logic;

begin
   
   Y_reg_28_inst : DLH_X1 port map( G => n4, D => N223, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n4, D => N222, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n4, D => N221, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n4, D => N220, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n4, D => N219, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n4, D => N218, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n4, D => N217, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n4, D => N216, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N215, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N214, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N213, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N212, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N211, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N210, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N209, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N208, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N207, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N206, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N205, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N204, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N203, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N202, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N201, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N200, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N199, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N198, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N197, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N196, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N195, Q => Y(0));
   n4 <= '1';
   U3 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n137, ZN => n16);
   U4 : OR4_X1 port map( A1 => n9, A2 => n7, A3 => n8, A4 => n134, ZN => n14);
   U5 : INV_X2 port map( A => n14, ZN => n1);
   U6 : OR3_X1 port map( A1 => n135, A2 => SEL(1), A3 => n137, ZN => n19);
   U7 : INV_X2 port map( A => n19, ZN => n2);
   U8 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n135, ZN => n21);
   U9 : INV_X2 port map( A => n21, ZN => n3);
   U10 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n136, ZN => n18);
   U11 : INV_X2 port map( A => n18, ZN => n5);
   U12 : OR3_X1 port map( A1 => n137, A2 => n135, A3 => n136, ZN => n20);
   U13 : INV_X2 port map( A => n20, ZN => n6);
   U14 : OR3_X1 port map( A1 => n137, A2 => SEL(2), A3 => n136, ZN => n17);
   U15 : INV_X2 port map( A => n17, ZN => n7);
   U16 : OR3_X1 port map( A1 => n135, A2 => SEL(0), A3 => n136, ZN => n15);
   U17 : INV_X2 port map( A => n15, ZN => n8);
   U18 : CLKBUF_X2 port map( A => n16, Z => n9);
   U19 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           N223);
   U20 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(174), B2 =>
                           n8, ZN => n13);
   U21 : AOI22_X1 port map( A1 => inputs(29), A2 => n9, B1 => inputs(87), B2 =>
                           n7, ZN => n12);
   U22 : AOI22_X1 port map( A1 => inputs(58), A2 => n5, B1 => inputs(145), B2 
                           => n2, ZN => n11);
   U23 : AOI22_X1 port map( A1 => inputs(203), A2 => n6, B1 => inputs(116), B2 
                           => n3, ZN => n10);
   U24 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           N222);
   U25 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(175), B2 =>
                           n8, ZN => n25);
   U26 : AOI22_X1 port map( A1 => inputs(30), A2 => n9, B1 => inputs(88), B2 =>
                           n7, ZN => n24);
   U27 : AOI22_X1 port map( A1 => inputs(59), A2 => n5, B1 => inputs(146), B2 
                           => n2, ZN => n23);
   U28 : AOI22_X1 port map( A1 => inputs(204), A2 => n6, B1 => inputs(117), B2 
                           => n3, ZN => n22);
   U29 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n28, A4 => n29, ZN => 
                           N221);
   U30 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(176), B2 =>
                           n8, ZN => n29);
   U31 : AOI22_X1 port map( A1 => inputs(31), A2 => n9, B1 => inputs(89), B2 =>
                           n7, ZN => n28);
   U32 : AOI22_X1 port map( A1 => inputs(60), A2 => n5, B1 => inputs(147), B2 
                           => n2, ZN => n27);
   U33 : AOI22_X1 port map( A1 => inputs(205), A2 => n6, B1 => inputs(118), B2 
                           => n3, ZN => n26);
   U34 : NAND4_X1 port map( A1 => n30, A2 => n31, A3 => n32, A4 => n33, ZN => 
                           N220);
   U35 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(177), B2 =>
                           n8, ZN => n33);
   U36 : AOI22_X1 port map( A1 => inputs(32), A2 => n9, B1 => inputs(90), B2 =>
                           n7, ZN => n32);
   U37 : AOI22_X1 port map( A1 => inputs(61), A2 => n5, B1 => inputs(148), B2 
                           => n2, ZN => n31);
   U38 : AOI22_X1 port map( A1 => inputs(206), A2 => n6, B1 => inputs(119), B2 
                           => n3, ZN => n30);
   U39 : NAND4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           N219);
   U40 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(178), B2 =>
                           n8, ZN => n37);
   U41 : AOI22_X1 port map( A1 => inputs(33), A2 => n9, B1 => inputs(91), B2 =>
                           n7, ZN => n36);
   U42 : AOI22_X1 port map( A1 => inputs(62), A2 => n5, B1 => inputs(149), B2 
                           => n2, ZN => n35);
   U43 : AOI22_X1 port map( A1 => inputs(207), A2 => n6, B1 => inputs(120), B2 
                           => n3, ZN => n34);
   U44 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           N218);
   U45 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(179), B2 =>
                           n8, ZN => n41);
   U46 : AOI22_X1 port map( A1 => inputs(34), A2 => n9, B1 => inputs(92), B2 =>
                           n7, ZN => n40);
   U47 : AOI22_X1 port map( A1 => inputs(63), A2 => n5, B1 => inputs(150), B2 
                           => n2, ZN => n39);
   U48 : AOI22_X1 port map( A1 => inputs(208), A2 => n6, B1 => inputs(121), B2 
                           => n3, ZN => n38);
   U49 : NAND4_X1 port map( A1 => n42, A2 => n43, A3 => n44, A4 => n45, ZN => 
                           N217);
   U50 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(180), B2 =>
                           n8, ZN => n45);
   U51 : AOI22_X1 port map( A1 => inputs(35), A2 => n9, B1 => inputs(93), B2 =>
                           n7, ZN => n44);
   U52 : AOI22_X1 port map( A1 => inputs(64), A2 => n5, B1 => inputs(151), B2 
                           => n2, ZN => n43);
   U53 : AOI22_X1 port map( A1 => inputs(209), A2 => n6, B1 => inputs(122), B2 
                           => n3, ZN => n42);
   U54 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           N216);
   U55 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(181), B2 =>
                           n8, ZN => n49);
   U56 : AOI22_X1 port map( A1 => inputs(36), A2 => n9, B1 => inputs(94), B2 =>
                           n7, ZN => n48);
   U57 : AOI22_X1 port map( A1 => inputs(65), A2 => n5, B1 => inputs(152), B2 
                           => n2, ZN => n47);
   U58 : AOI22_X1 port map( A1 => inputs(210), A2 => n6, B1 => inputs(123), B2 
                           => n3, ZN => n46);
   U59 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           N215);
   U60 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(182), B2 =>
                           n8, ZN => n53);
   U61 : AOI22_X1 port map( A1 => inputs(37), A2 => n9, B1 => inputs(95), B2 =>
                           n7, ZN => n52);
   U62 : AOI22_X1 port map( A1 => inputs(66), A2 => n5, B1 => inputs(153), B2 
                           => n2, ZN => n51);
   U63 : AOI22_X1 port map( A1 => inputs(211), A2 => n6, B1 => inputs(124), B2 
                           => n3, ZN => n50);
   U64 : NAND4_X1 port map( A1 => n54, A2 => n55, A3 => n56, A4 => n57, ZN => 
                           N214);
   U65 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(183), B2 =>
                           n8, ZN => n57);
   U66 : AOI22_X1 port map( A1 => inputs(38), A2 => n9, B1 => inputs(96), B2 =>
                           n7, ZN => n56);
   U67 : AOI22_X1 port map( A1 => inputs(67), A2 => n5, B1 => inputs(154), B2 
                           => n2, ZN => n55);
   U68 : AOI22_X1 port map( A1 => inputs(212), A2 => n6, B1 => inputs(125), B2 
                           => n3, ZN => n54);
   U69 : NAND4_X1 port map( A1 => n58, A2 => n59, A3 => n60, A4 => n61, ZN => 
                           N213);
   U70 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(184), B2 
                           => n8, ZN => n61);
   U71 : AOI22_X1 port map( A1 => inputs(39), A2 => n9, B1 => inputs(97), B2 =>
                           n7, ZN => n60);
   U72 : AOI22_X1 port map( A1 => inputs(68), A2 => n5, B1 => inputs(155), B2 
                           => n2, ZN => n59);
   U73 : AOI22_X1 port map( A1 => inputs(213), A2 => n6, B1 => inputs(126), B2 
                           => n3, ZN => n58);
   U74 : NAND4_X1 port map( A1 => n62, A2 => n63, A3 => n64, A4 => n65, ZN => 
                           N212);
   U75 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(185), B2 
                           => n8, ZN => n65);
   U76 : AOI22_X1 port map( A1 => inputs(40), A2 => n9, B1 => inputs(98), B2 =>
                           n7, ZN => n64);
   U77 : AOI22_X1 port map( A1 => inputs(69), A2 => n5, B1 => inputs(156), B2 
                           => n2, ZN => n63);
   U78 : AOI22_X1 port map( A1 => inputs(214), A2 => n6, B1 => inputs(127), B2 
                           => n3, ZN => n62);
   U79 : NAND4_X1 port map( A1 => n66, A2 => n67, A3 => n68, A4 => n69, ZN => 
                           N211);
   U80 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(186), B2 
                           => n8, ZN => n69);
   U81 : AOI22_X1 port map( A1 => inputs(41), A2 => n9, B1 => inputs(99), B2 =>
                           n7, ZN => n68);
   U82 : AOI22_X1 port map( A1 => inputs(70), A2 => n5, B1 => inputs(157), B2 
                           => n2, ZN => n67);
   U83 : AOI22_X1 port map( A1 => inputs(215), A2 => n6, B1 => inputs(128), B2 
                           => n3, ZN => n66);
   U84 : NAND4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           N210);
   U85 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(187), B2 
                           => n8, ZN => n73);
   U86 : AOI22_X1 port map( A1 => inputs(42), A2 => n9, B1 => inputs(100), B2 
                           => n7, ZN => n72);
   U87 : AOI22_X1 port map( A1 => inputs(71), A2 => n5, B1 => inputs(158), B2 
                           => n2, ZN => n71);
   U88 : AOI22_X1 port map( A1 => inputs(216), A2 => n6, B1 => inputs(129), B2 
                           => n3, ZN => n70);
   U89 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           N209);
   U90 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(188), B2 
                           => n8, ZN => n77);
   U91 : AOI22_X1 port map( A1 => inputs(43), A2 => n9, B1 => inputs(101), B2 
                           => n7, ZN => n76);
   U92 : AOI22_X1 port map( A1 => inputs(72), A2 => n5, B1 => inputs(159), B2 
                           => n2, ZN => n75);
   U93 : AOI22_X1 port map( A1 => inputs(217), A2 => n6, B1 => inputs(130), B2 
                           => n3, ZN => n74);
   U94 : NAND4_X1 port map( A1 => n78, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           N208);
   U95 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(189), B2 
                           => n8, ZN => n81);
   U96 : AOI22_X1 port map( A1 => inputs(44), A2 => n9, B1 => inputs(102), B2 
                           => n7, ZN => n80);
   U97 : AOI22_X1 port map( A1 => inputs(73), A2 => n5, B1 => inputs(160), B2 
                           => n2, ZN => n79);
   U98 : AOI22_X1 port map( A1 => inputs(218), A2 => n6, B1 => inputs(131), B2 
                           => n3, ZN => n78);
   U99 : NAND4_X1 port map( A1 => n82, A2 => n83, A3 => n84, A4 => n85, ZN => 
                           N207);
   U100 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(190), B2 
                           => n8, ZN => n85);
   U101 : AOI22_X1 port map( A1 => inputs(45), A2 => n9, B1 => inputs(103), B2 
                           => n7, ZN => n84);
   U102 : AOI22_X1 port map( A1 => inputs(74), A2 => n5, B1 => inputs(161), B2 
                           => n2, ZN => n83);
   U103 : AOI22_X1 port map( A1 => inputs(219), A2 => n6, B1 => inputs(132), B2
                           => n3, ZN => n82);
   U104 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           N206);
   U105 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(191), B2 
                           => n8, ZN => n89);
   U106 : AOI22_X1 port map( A1 => inputs(46), A2 => n9, B1 => inputs(104), B2 
                           => n7, ZN => n88);
   U107 : AOI22_X1 port map( A1 => inputs(75), A2 => n5, B1 => inputs(162), B2 
                           => n2, ZN => n87);
   U108 : AOI22_X1 port map( A1 => inputs(220), A2 => n6, B1 => inputs(133), B2
                           => n3, ZN => n86);
   U109 : NAND4_X1 port map( A1 => n90, A2 => n91, A3 => n92, A4 => n93, ZN => 
                           N205);
   U110 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(192), B2 
                           => n8, ZN => n93);
   U111 : AOI22_X1 port map( A1 => inputs(47), A2 => n9, B1 => inputs(105), B2 
                           => n7, ZN => n92);
   U112 : AOI22_X1 port map( A1 => inputs(76), A2 => n5, B1 => inputs(163), B2 
                           => n2, ZN => n91);
   U113 : AOI22_X1 port map( A1 => inputs(221), A2 => n6, B1 => inputs(134), B2
                           => n3, ZN => n90);
   U114 : NAND4_X1 port map( A1 => n94, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           N204);
   U115 : AOI22_X1 port map( A1 => inputs(19), A2 => n1, B1 => inputs(193), B2 
                           => n8, ZN => n97);
   U116 : AOI22_X1 port map( A1 => inputs(48), A2 => n9, B1 => inputs(106), B2 
                           => n7, ZN => n96);
   U117 : AOI22_X1 port map( A1 => inputs(77), A2 => n5, B1 => inputs(164), B2 
                           => n2, ZN => n95);
   U118 : AOI22_X1 port map( A1 => inputs(222), A2 => n6, B1 => inputs(135), B2
                           => n3, ZN => n94);
   U119 : NAND4_X1 port map( A1 => n98, A2 => n99, A3 => n100, A4 => n101, ZN 
                           => N203);
   U120 : AOI22_X1 port map( A1 => inputs(20), A2 => n1, B1 => inputs(194), B2 
                           => n8, ZN => n101);
   U121 : AOI22_X1 port map( A1 => inputs(49), A2 => n9, B1 => inputs(107), B2 
                           => n7, ZN => n100);
   U122 : AOI22_X1 port map( A1 => inputs(78), A2 => n5, B1 => inputs(165), B2 
                           => n2, ZN => n99);
   U123 : AOI22_X1 port map( A1 => inputs(223), A2 => n6, B1 => inputs(136), B2
                           => n3, ZN => n98);
   U124 : NAND4_X1 port map( A1 => n102, A2 => n103, A3 => n104, A4 => n105, ZN
                           => N202);
   U125 : AOI22_X1 port map( A1 => inputs(21), A2 => n1, B1 => inputs(195), B2 
                           => n8, ZN => n105);
   U126 : AOI22_X1 port map( A1 => inputs(50), A2 => n9, B1 => inputs(108), B2 
                           => n7, ZN => n104);
   U127 : AOI22_X1 port map( A1 => inputs(79), A2 => n5, B1 => inputs(166), B2 
                           => n2, ZN => n103);
   U128 : AOI22_X1 port map( A1 => inputs(224), A2 => n6, B1 => inputs(137), B2
                           => n3, ZN => n102);
   U129 : NAND4_X1 port map( A1 => n106, A2 => n107, A3 => n108, A4 => n109, ZN
                           => N201);
   U130 : AOI22_X1 port map( A1 => inputs(22), A2 => n1, B1 => inputs(196), B2 
                           => n8, ZN => n109);
   U131 : AOI22_X1 port map( A1 => inputs(51), A2 => n9, B1 => inputs(109), B2 
                           => n7, ZN => n108);
   U132 : AOI22_X1 port map( A1 => inputs(80), A2 => n5, B1 => inputs(167), B2 
                           => n2, ZN => n107);
   U133 : AOI22_X1 port map( A1 => inputs(225), A2 => n6, B1 => inputs(138), B2
                           => n3, ZN => n106);
   U134 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN
                           => N200);
   U135 : AOI22_X1 port map( A1 => inputs(23), A2 => n1, B1 => inputs(197), B2 
                           => n8, ZN => n113);
   U136 : AOI22_X1 port map( A1 => inputs(52), A2 => n9, B1 => inputs(110), B2 
                           => n7, ZN => n112);
   U137 : AOI22_X1 port map( A1 => inputs(81), A2 => n5, B1 => inputs(168), B2 
                           => n2, ZN => n111);
   U138 : AOI22_X1 port map( A1 => inputs(226), A2 => n6, B1 => inputs(139), B2
                           => n3, ZN => n110);
   U139 : NAND4_X1 port map( A1 => n114, A2 => n115, A3 => n116, A4 => n117, ZN
                           => N199);
   U140 : AOI22_X1 port map( A1 => inputs(24), A2 => n1, B1 => inputs(198), B2 
                           => n8, ZN => n117);
   U141 : AOI22_X1 port map( A1 => inputs(53), A2 => n9, B1 => inputs(111), B2 
                           => n7, ZN => n116);
   U142 : AOI22_X1 port map( A1 => inputs(82), A2 => n5, B1 => inputs(169), B2 
                           => n2, ZN => n115);
   U143 : AOI22_X1 port map( A1 => inputs(227), A2 => n6, B1 => inputs(140), B2
                           => n3, ZN => n114);
   U144 : NAND4_X1 port map( A1 => n118, A2 => n119, A3 => n120, A4 => n121, ZN
                           => N198);
   U145 : AOI22_X1 port map( A1 => inputs(25), A2 => n1, B1 => inputs(199), B2 
                           => n8, ZN => n121);
   U146 : AOI22_X1 port map( A1 => inputs(54), A2 => n9, B1 => inputs(112), B2 
                           => n7, ZN => n120);
   U147 : AOI22_X1 port map( A1 => inputs(83), A2 => n5, B1 => inputs(170), B2 
                           => n2, ZN => n119);
   U148 : AOI22_X1 port map( A1 => inputs(228), A2 => n6, B1 => inputs(141), B2
                           => n3, ZN => n118);
   U149 : NAND4_X1 port map( A1 => n122, A2 => n123, A3 => n124, A4 => n125, ZN
                           => N197);
   U150 : AOI22_X1 port map( A1 => inputs(26), A2 => n1, B1 => inputs(200), B2 
                           => n8, ZN => n125);
   U151 : AOI22_X1 port map( A1 => inputs(55), A2 => n9, B1 => inputs(113), B2 
                           => n7, ZN => n124);
   U152 : AOI22_X1 port map( A1 => inputs(84), A2 => n5, B1 => inputs(171), B2 
                           => n2, ZN => n123);
   U153 : AOI22_X1 port map( A1 => inputs(229), A2 => n6, B1 => inputs(142), B2
                           => n3, ZN => n122);
   U154 : NAND4_X1 port map( A1 => n126, A2 => n127, A3 => n128, A4 => n129, ZN
                           => N196);
   U155 : AOI22_X1 port map( A1 => inputs(27), A2 => n1, B1 => inputs(201), B2 
                           => n8, ZN => n129);
   U156 : AOI22_X1 port map( A1 => inputs(56), A2 => n9, B1 => inputs(114), B2 
                           => n7, ZN => n128);
   U157 : AOI22_X1 port map( A1 => inputs(85), A2 => n5, B1 => inputs(172), B2 
                           => n2, ZN => n127);
   U158 : AOI22_X1 port map( A1 => inputs(230), A2 => n6, B1 => inputs(143), B2
                           => n3, ZN => n126);
   U159 : NAND4_X1 port map( A1 => n130, A2 => n131, A3 => n132, A4 => n133, ZN
                           => N195);
   U161 : AOI22_X1 port map( A1 => inputs(28), A2 => n1, B1 => inputs(202), B2 
                           => n8, ZN => n133);
   U162 : OR4_X1 port map( A1 => n3, A2 => n6, A3 => n2, A4 => n5, ZN => n134);
   U163 : AOI22_X1 port map( A1 => inputs(57), A2 => n9, B1 => inputs(115), B2 
                           => n7, ZN => n132);
   U164 : AOI22_X1 port map( A1 => inputs(86), A2 => n5, B1 => inputs(173), B2 
                           => n2, ZN => n131);
   U165 : AOI22_X1 port map( A1 => inputs(231), A2 => n6, B1 => inputs(144), B2
                           => n3, ZN => n130);
   U166 : INV_X1 port map( A => SEL(1), ZN => n136);
   U167 : INV_X1 port map( A => SEL(2), ZN => n135);
   U168 : INV_X1 port map( A => SEL(0), ZN => n137);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT27 is

   port( a, b : in std_logic_vector (26 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (27 downto 0));

end adder_NBIT27;

architecture SYN_beh of adder_NBIT27 is

   component adder_NBIT27_DW01_add_0
      port( A, B : in std_logic_vector (27 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (27 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3351 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT27_DW01_add_0 port map( A(27) => a(26), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), B(27) => b(26), B(26) => b(26), 
                           B(25) => b(25), B(24) => b(24), B(23) => b(23), 
                           B(22) => b(22), B(21) => b(21), B(20) => b(20), 
                           B(19) => b(19), B(18) => b(18), B(17) => b(17), 
                           B(16) => b(16), B(15) => b(15), B(14) => b(14), 
                           B(13) => b(13), B(12) => b(12), B(11) => b(11), 
                           B(10) => b(10), B(9) => b(9), B(8) => b(8), B(7) => 
                           b(7), B(6) => b(6), B(5) => b(5), B(4) => b(4), B(3)
                           => b(3), B(2) => b(2), B(1) => b(1), B(0) => b(0), 
                           CI => cin, SUM(27) => s(27), SUM(26) => s(26), 
                           SUM(25) => s(25), SUM(24) => s(24), SUM(23) => s(23)
                           , SUM(22) => s(22), SUM(21) => s(21), SUM(20) => 
                           s(20), SUM(19) => s(19), SUM(18) => s(18), SUM(17) 
                           => s(17), SUM(16) => s(16), SUM(15) => s(15), 
                           SUM(14) => s(14), SUM(13) => s(13), SUM(12) => s(12)
                           , SUM(11) => s(11), SUM(10) => s(10), SUM(9) => s(9)
                           , SUM(8) => s(8), SUM(7) => s(7), SUM(6) => s(6), 
                           SUM(5) => s(5), SUM(4) => s(4), SUM(3) => s(3), 
                           SUM(2) => s(2), SUM(1) => s(1), SUM(0) => s(0), CO 
                           => n_3351);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N27_Z3 is

   port( inputs : in std_logic_vector (0 to 215);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (26 downto 0));

end MUX_zbit_nbit_N27_Z3;

architecture SYN_beh of MUX_zbit_nbit_N27_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, 
      N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, 
      N206, N207, N208, N209, n4, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129 : std_logic;

begin
   
   Y_reg_26_inst : DLH_X1 port map( G => n4, D => N209, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n4, D => N208, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n4, D => N207, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n4, D => N206, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n4, D => N205, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n4, D => N204, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N203, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N202, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N201, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N200, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N199, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N198, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N197, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N196, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N195, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N194, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N193, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N192, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N191, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N190, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N189, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N188, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N187, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N186, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N185, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N184, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N183, Q => Y(0));
   n4 <= '1';
   U3 : OR4_X1 port map( A1 => n9, A2 => n7, A3 => n8, A4 => n126, ZN => n14);
   U4 : INV_X2 port map( A => n14, ZN => n1);
   U5 : OR3_X1 port map( A1 => n127, A2 => SEL(1), A3 => n129, ZN => n19);
   U6 : INV_X2 port map( A => n19, ZN => n2);
   U7 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n127, ZN => n21);
   U8 : INV_X2 port map( A => n21, ZN => n3);
   U9 : OR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n128, ZN => n18);
   U10 : INV_X2 port map( A => n18, ZN => n5);
   U11 : OR3_X1 port map( A1 => n129, A2 => n127, A3 => n128, ZN => n20);
   U12 : INV_X2 port map( A => n20, ZN => n6);
   U13 : OR3_X1 port map( A1 => n129, A2 => SEL(2), A3 => n128, ZN => n17);
   U14 : INV_X2 port map( A => n17, ZN => n7);
   U15 : OR3_X1 port map( A1 => n127, A2 => SEL(0), A3 => n128, ZN => n15);
   U16 : INV_X2 port map( A => n15, ZN => n8);
   U17 : OR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n129, ZN => n16);
   U18 : INV_X2 port map( A => n16, ZN => n9);
   U19 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           N209);
   U20 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(162), B2 =>
                           n8, ZN => n13);
   U21 : AOI22_X1 port map( A1 => inputs(27), A2 => n9, B1 => inputs(81), B2 =>
                           n7, ZN => n12);
   U22 : AOI22_X1 port map( A1 => inputs(54), A2 => n5, B1 => inputs(135), B2 
                           => n2, ZN => n11);
   U23 : AOI22_X1 port map( A1 => inputs(189), A2 => n6, B1 => inputs(108), B2 
                           => n3, ZN => n10);
   U24 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           N208);
   U25 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(163), B2 =>
                           n8, ZN => n25);
   U26 : AOI22_X1 port map( A1 => inputs(28), A2 => n9, B1 => inputs(82), B2 =>
                           n7, ZN => n24);
   U27 : AOI22_X1 port map( A1 => inputs(55), A2 => n5, B1 => inputs(136), B2 
                           => n2, ZN => n23);
   U28 : AOI22_X1 port map( A1 => inputs(190), A2 => n6, B1 => inputs(109), B2 
                           => n3, ZN => n22);
   U29 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n28, A4 => n29, ZN => 
                           N207);
   U30 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(164), B2 =>
                           n8, ZN => n29);
   U31 : AOI22_X1 port map( A1 => inputs(29), A2 => n9, B1 => inputs(83), B2 =>
                           n7, ZN => n28);
   U32 : AOI22_X1 port map( A1 => inputs(56), A2 => n5, B1 => inputs(137), B2 
                           => n2, ZN => n27);
   U33 : AOI22_X1 port map( A1 => inputs(191), A2 => n6, B1 => inputs(110), B2 
                           => n3, ZN => n26);
   U34 : NAND4_X1 port map( A1 => n30, A2 => n31, A3 => n32, A4 => n33, ZN => 
                           N206);
   U35 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(165), B2 =>
                           n8, ZN => n33);
   U36 : AOI22_X1 port map( A1 => inputs(30), A2 => n9, B1 => inputs(84), B2 =>
                           n7, ZN => n32);
   U37 : AOI22_X1 port map( A1 => inputs(57), A2 => n5, B1 => inputs(138), B2 
                           => n2, ZN => n31);
   U38 : AOI22_X1 port map( A1 => inputs(192), A2 => n6, B1 => inputs(111), B2 
                           => n3, ZN => n30);
   U39 : NAND4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           N205);
   U40 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(166), B2 =>
                           n8, ZN => n37);
   U41 : AOI22_X1 port map( A1 => inputs(31), A2 => n9, B1 => inputs(85), B2 =>
                           n7, ZN => n36);
   U42 : AOI22_X1 port map( A1 => inputs(58), A2 => n5, B1 => inputs(139), B2 
                           => n2, ZN => n35);
   U43 : AOI22_X1 port map( A1 => inputs(193), A2 => n6, B1 => inputs(112), B2 
                           => n3, ZN => n34);
   U44 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           N204);
   U45 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(167), B2 =>
                           n8, ZN => n41);
   U46 : AOI22_X1 port map( A1 => inputs(32), A2 => n9, B1 => inputs(86), B2 =>
                           n7, ZN => n40);
   U47 : AOI22_X1 port map( A1 => inputs(59), A2 => n5, B1 => inputs(140), B2 
                           => n2, ZN => n39);
   U48 : AOI22_X1 port map( A1 => inputs(194), A2 => n6, B1 => inputs(113), B2 
                           => n3, ZN => n38);
   U49 : NAND4_X1 port map( A1 => n42, A2 => n43, A3 => n44, A4 => n45, ZN => 
                           N203);
   U50 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(168), B2 =>
                           n8, ZN => n45);
   U51 : AOI22_X1 port map( A1 => inputs(33), A2 => n9, B1 => inputs(87), B2 =>
                           n7, ZN => n44);
   U52 : AOI22_X1 port map( A1 => inputs(60), A2 => n5, B1 => inputs(141), B2 
                           => n2, ZN => n43);
   U53 : AOI22_X1 port map( A1 => inputs(195), A2 => n6, B1 => inputs(114), B2 
                           => n3, ZN => n42);
   U54 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           N202);
   U55 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(169), B2 =>
                           n8, ZN => n49);
   U56 : AOI22_X1 port map( A1 => inputs(34), A2 => n9, B1 => inputs(88), B2 =>
                           n7, ZN => n48);
   U57 : AOI22_X1 port map( A1 => inputs(61), A2 => n5, B1 => inputs(142), B2 
                           => n2, ZN => n47);
   U58 : AOI22_X1 port map( A1 => inputs(196), A2 => n6, B1 => inputs(115), B2 
                           => n3, ZN => n46);
   U59 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           N201);
   U60 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(170), B2 =>
                           n8, ZN => n53);
   U61 : AOI22_X1 port map( A1 => inputs(35), A2 => n9, B1 => inputs(89), B2 =>
                           n7, ZN => n52);
   U62 : AOI22_X1 port map( A1 => inputs(62), A2 => n5, B1 => inputs(143), B2 
                           => n2, ZN => n51);
   U63 : AOI22_X1 port map( A1 => inputs(197), A2 => n6, B1 => inputs(116), B2 
                           => n3, ZN => n50);
   U64 : NAND4_X1 port map( A1 => n54, A2 => n55, A3 => n56, A4 => n57, ZN => 
                           N200);
   U65 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(171), B2 =>
                           n8, ZN => n57);
   U66 : AOI22_X1 port map( A1 => inputs(36), A2 => n9, B1 => inputs(90), B2 =>
                           n7, ZN => n56);
   U67 : AOI22_X1 port map( A1 => inputs(63), A2 => n5, B1 => inputs(144), B2 
                           => n2, ZN => n55);
   U68 : AOI22_X1 port map( A1 => inputs(198), A2 => n6, B1 => inputs(117), B2 
                           => n3, ZN => n54);
   U69 : NAND4_X1 port map( A1 => n58, A2 => n59, A3 => n60, A4 => n61, ZN => 
                           N199);
   U70 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(172), B2 
                           => n8, ZN => n61);
   U71 : AOI22_X1 port map( A1 => inputs(37), A2 => n9, B1 => inputs(91), B2 =>
                           n7, ZN => n60);
   U72 : AOI22_X1 port map( A1 => inputs(64), A2 => n5, B1 => inputs(145), B2 
                           => n2, ZN => n59);
   U73 : AOI22_X1 port map( A1 => inputs(199), A2 => n6, B1 => inputs(118), B2 
                           => n3, ZN => n58);
   U74 : NAND4_X1 port map( A1 => n62, A2 => n63, A3 => n64, A4 => n65, ZN => 
                           N198);
   U75 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(173), B2 
                           => n8, ZN => n65);
   U76 : AOI22_X1 port map( A1 => inputs(38), A2 => n9, B1 => inputs(92), B2 =>
                           n7, ZN => n64);
   U77 : AOI22_X1 port map( A1 => inputs(65), A2 => n5, B1 => inputs(146), B2 
                           => n2, ZN => n63);
   U78 : AOI22_X1 port map( A1 => inputs(200), A2 => n6, B1 => inputs(119), B2 
                           => n3, ZN => n62);
   U79 : NAND4_X1 port map( A1 => n66, A2 => n67, A3 => n68, A4 => n69, ZN => 
                           N197);
   U80 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(174), B2 
                           => n8, ZN => n69);
   U81 : AOI22_X1 port map( A1 => inputs(39), A2 => n9, B1 => inputs(93), B2 =>
                           n7, ZN => n68);
   U82 : AOI22_X1 port map( A1 => inputs(66), A2 => n5, B1 => inputs(147), B2 
                           => n2, ZN => n67);
   U83 : AOI22_X1 port map( A1 => inputs(201), A2 => n6, B1 => inputs(120), B2 
                           => n3, ZN => n66);
   U84 : NAND4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           N196);
   U85 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(175), B2 
                           => n8, ZN => n73);
   U86 : AOI22_X1 port map( A1 => inputs(40), A2 => n9, B1 => inputs(94), B2 =>
                           n7, ZN => n72);
   U87 : AOI22_X1 port map( A1 => inputs(67), A2 => n5, B1 => inputs(148), B2 
                           => n2, ZN => n71);
   U88 : AOI22_X1 port map( A1 => inputs(202), A2 => n6, B1 => inputs(121), B2 
                           => n3, ZN => n70);
   U89 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           N195);
   U90 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(176), B2 
                           => n8, ZN => n77);
   U91 : AOI22_X1 port map( A1 => inputs(41), A2 => n9, B1 => inputs(95), B2 =>
                           n7, ZN => n76);
   U92 : AOI22_X1 port map( A1 => inputs(68), A2 => n5, B1 => inputs(149), B2 
                           => n2, ZN => n75);
   U93 : AOI22_X1 port map( A1 => inputs(203), A2 => n6, B1 => inputs(122), B2 
                           => n3, ZN => n74);
   U94 : NAND4_X1 port map( A1 => n78, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           N194);
   U95 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(177), B2 
                           => n8, ZN => n81);
   U96 : AOI22_X1 port map( A1 => inputs(42), A2 => n9, B1 => inputs(96), B2 =>
                           n7, ZN => n80);
   U97 : AOI22_X1 port map( A1 => inputs(69), A2 => n5, B1 => inputs(150), B2 
                           => n2, ZN => n79);
   U98 : AOI22_X1 port map( A1 => inputs(204), A2 => n6, B1 => inputs(123), B2 
                           => n3, ZN => n78);
   U99 : NAND4_X1 port map( A1 => n82, A2 => n83, A3 => n84, A4 => n85, ZN => 
                           N193);
   U100 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(178), B2 
                           => n8, ZN => n85);
   U101 : AOI22_X1 port map( A1 => inputs(43), A2 => n9, B1 => inputs(97), B2 
                           => n7, ZN => n84);
   U102 : AOI22_X1 port map( A1 => inputs(70), A2 => n5, B1 => inputs(151), B2 
                           => n2, ZN => n83);
   U103 : AOI22_X1 port map( A1 => inputs(205), A2 => n6, B1 => inputs(124), B2
                           => n3, ZN => n82);
   U104 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           N192);
   U105 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(179), B2 
                           => n8, ZN => n89);
   U106 : AOI22_X1 port map( A1 => inputs(44), A2 => n9, B1 => inputs(98), B2 
                           => n7, ZN => n88);
   U107 : AOI22_X1 port map( A1 => inputs(71), A2 => n5, B1 => inputs(152), B2 
                           => n2, ZN => n87);
   U108 : AOI22_X1 port map( A1 => inputs(206), A2 => n6, B1 => inputs(125), B2
                           => n3, ZN => n86);
   U109 : NAND4_X1 port map( A1 => n90, A2 => n91, A3 => n92, A4 => n93, ZN => 
                           N191);
   U110 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(180), B2 
                           => n8, ZN => n93);
   U111 : AOI22_X1 port map( A1 => inputs(45), A2 => n9, B1 => inputs(99), B2 
                           => n7, ZN => n92);
   U112 : AOI22_X1 port map( A1 => inputs(72), A2 => n5, B1 => inputs(153), B2 
                           => n2, ZN => n91);
   U113 : AOI22_X1 port map( A1 => inputs(207), A2 => n6, B1 => inputs(126), B2
                           => n3, ZN => n90);
   U114 : NAND4_X1 port map( A1 => n94, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           N190);
   U115 : AOI22_X1 port map( A1 => inputs(19), A2 => n1, B1 => inputs(181), B2 
                           => n8, ZN => n97);
   U116 : AOI22_X1 port map( A1 => inputs(46), A2 => n9, B1 => inputs(100), B2 
                           => n7, ZN => n96);
   U117 : AOI22_X1 port map( A1 => inputs(73), A2 => n5, B1 => inputs(154), B2 
                           => n2, ZN => n95);
   U118 : AOI22_X1 port map( A1 => inputs(208), A2 => n6, B1 => inputs(127), B2
                           => n3, ZN => n94);
   U119 : NAND4_X1 port map( A1 => n98, A2 => n99, A3 => n100, A4 => n101, ZN 
                           => N189);
   U120 : AOI22_X1 port map( A1 => inputs(20), A2 => n1, B1 => inputs(182), B2 
                           => n8, ZN => n101);
   U121 : AOI22_X1 port map( A1 => inputs(47), A2 => n9, B1 => inputs(101), B2 
                           => n7, ZN => n100);
   U122 : AOI22_X1 port map( A1 => inputs(74), A2 => n5, B1 => inputs(155), B2 
                           => n2, ZN => n99);
   U123 : AOI22_X1 port map( A1 => inputs(209), A2 => n6, B1 => inputs(128), B2
                           => n3, ZN => n98);
   U124 : NAND4_X1 port map( A1 => n102, A2 => n103, A3 => n104, A4 => n105, ZN
                           => N188);
   U125 : AOI22_X1 port map( A1 => inputs(21), A2 => n1, B1 => inputs(183), B2 
                           => n8, ZN => n105);
   U126 : AOI22_X1 port map( A1 => inputs(48), A2 => n9, B1 => inputs(102), B2 
                           => n7, ZN => n104);
   U127 : AOI22_X1 port map( A1 => inputs(75), A2 => n5, B1 => inputs(156), B2 
                           => n2, ZN => n103);
   U128 : AOI22_X1 port map( A1 => inputs(210), A2 => n6, B1 => inputs(129), B2
                           => n3, ZN => n102);
   U129 : NAND4_X1 port map( A1 => n106, A2 => n107, A3 => n108, A4 => n109, ZN
                           => N187);
   U130 : AOI22_X1 port map( A1 => inputs(22), A2 => n1, B1 => inputs(184), B2 
                           => n8, ZN => n109);
   U131 : AOI22_X1 port map( A1 => inputs(49), A2 => n9, B1 => inputs(103), B2 
                           => n7, ZN => n108);
   U132 : AOI22_X1 port map( A1 => inputs(76), A2 => n5, B1 => inputs(157), B2 
                           => n2, ZN => n107);
   U133 : AOI22_X1 port map( A1 => inputs(211), A2 => n6, B1 => inputs(130), B2
                           => n3, ZN => n106);
   U134 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN
                           => N186);
   U135 : AOI22_X1 port map( A1 => inputs(23), A2 => n1, B1 => inputs(185), B2 
                           => n8, ZN => n113);
   U136 : AOI22_X1 port map( A1 => inputs(50), A2 => n9, B1 => inputs(104), B2 
                           => n7, ZN => n112);
   U137 : AOI22_X1 port map( A1 => inputs(77), A2 => n5, B1 => inputs(158), B2 
                           => n2, ZN => n111);
   U138 : AOI22_X1 port map( A1 => inputs(212), A2 => n6, B1 => inputs(131), B2
                           => n3, ZN => n110);
   U139 : NAND4_X1 port map( A1 => n114, A2 => n115, A3 => n116, A4 => n117, ZN
                           => N185);
   U140 : AOI22_X1 port map( A1 => inputs(24), A2 => n1, B1 => inputs(186), B2 
                           => n8, ZN => n117);
   U141 : AOI22_X1 port map( A1 => inputs(51), A2 => n9, B1 => inputs(105), B2 
                           => n7, ZN => n116);
   U142 : AOI22_X1 port map( A1 => inputs(78), A2 => n5, B1 => inputs(159), B2 
                           => n2, ZN => n115);
   U143 : AOI22_X1 port map( A1 => inputs(213), A2 => n6, B1 => inputs(132), B2
                           => n3, ZN => n114);
   U144 : NAND4_X1 port map( A1 => n118, A2 => n119, A3 => n120, A4 => n121, ZN
                           => N184);
   U145 : AOI22_X1 port map( A1 => inputs(25), A2 => n1, B1 => inputs(187), B2 
                           => n8, ZN => n121);
   U146 : AOI22_X1 port map( A1 => inputs(52), A2 => n9, B1 => inputs(106), B2 
                           => n7, ZN => n120);
   U147 : AOI22_X1 port map( A1 => inputs(79), A2 => n5, B1 => inputs(160), B2 
                           => n2, ZN => n119);
   U148 : AOI22_X1 port map( A1 => inputs(214), A2 => n6, B1 => inputs(133), B2
                           => n3, ZN => n118);
   U149 : NAND4_X1 port map( A1 => n122, A2 => n123, A3 => n124, A4 => n125, ZN
                           => N183);
   U151 : AOI22_X1 port map( A1 => inputs(26), A2 => n1, B1 => inputs(188), B2 
                           => n8, ZN => n125);
   U152 : OR4_X1 port map( A1 => n3, A2 => n6, A3 => n2, A4 => n5, ZN => n126);
   U153 : AOI22_X1 port map( A1 => inputs(53), A2 => n9, B1 => inputs(107), B2 
                           => n7, ZN => n124);
   U154 : AOI22_X1 port map( A1 => inputs(80), A2 => n5, B1 => inputs(161), B2 
                           => n2, ZN => n123);
   U155 : AOI22_X1 port map( A1 => inputs(215), A2 => n6, B1 => inputs(134), B2
                           => n3, ZN => n122);
   U156 : INV_X1 port map( A => SEL(1), ZN => n128);
   U157 : INV_X1 port map( A => SEL(2), ZN => n127);
   U158 : INV_X1 port map( A => SEL(0), ZN => n129);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT25 is

   port( a, b : in std_logic_vector (24 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (25 downto 0));

end adder_NBIT25;

architecture SYN_beh of adder_NBIT25 is

   component adder_NBIT25_DW01_add_0
      port( A, B : in std_logic_vector (25 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (25 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3352 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT25_DW01_add_0 port map( A(25) => a(24), 
                           A(24) => a(24), A(23) => a(23), A(22) => a(22), 
                           A(21) => a(21), A(20) => a(20), A(19) => a(19), 
                           A(18) => a(18), A(17) => a(17), A(16) => a(16), 
                           A(15) => a(15), A(14) => a(14), A(13) => a(13), 
                           A(12) => a(12), A(11) => a(11), A(10) => a(10), A(9)
                           => a(9), A(8) => a(8), A(7) => a(7), A(6) => a(6), 
                           A(5) => a(5), A(4) => a(4), A(3) => a(3), A(2) => 
                           a(2), A(1) => a(1), A(0) => a(0), B(25) => b(24), 
                           B(24) => b(24), B(23) => b(23), B(22) => b(22), 
                           B(21) => b(21), B(20) => b(20), B(19) => b(19), 
                           B(18) => b(18), B(17) => b(17), B(16) => b(16), 
                           B(15) => b(15), B(14) => b(14), B(13) => b(13), 
                           B(12) => b(12), B(11) => b(11), B(10) => b(10), B(9)
                           => b(9), B(8) => b(8), B(7) => b(7), B(6) => b(6), 
                           B(5) => b(5), B(4) => b(4), B(3) => b(3), B(2) => 
                           b(2), B(1) => b(1), B(0) => b(0), CI => cin, SUM(25)
                           => s(25), SUM(24) => s(24), SUM(23) => s(23), 
                           SUM(22) => s(22), SUM(21) => s(21), SUM(20) => s(20)
                           , SUM(19) => s(19), SUM(18) => s(18), SUM(17) => 
                           s(17), SUM(16) => s(16), SUM(15) => s(15), SUM(14) 
                           => s(14), SUM(13) => s(13), SUM(12) => s(12), 
                           SUM(11) => s(11), SUM(10) => s(10), SUM(9) => s(9), 
                           SUM(8) => s(8), SUM(7) => s(7), SUM(6) => s(6), 
                           SUM(5) => s(5), SUM(4) => s(4), SUM(3) => s(3), 
                           SUM(2) => s(2), SUM(1) => s(1), SUM(0) => s(0), CO 
                           => n_3352);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N25_Z3 is

   port( inputs : in std_logic_vector (0 to 199);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (24 downto 0));

end MUX_zbit_nbit_N25_Z3;

architecture SYN_beh of MUX_zbit_nbit_N25_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, 
      N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, 
      N194, N195, n4, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117 : std_logic;

begin
   
   Y_reg_24_inst : DLH_X1 port map( G => n4, D => N195, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n4, D => N194, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n4, D => N193, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n4, D => N192, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N191, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N190, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N189, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N188, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N187, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N186, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N185, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N184, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N183, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N182, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N181, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N180, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N179, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N178, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N177, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N176, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N175, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N174, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N173, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N172, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N171, Q => Y(0));
   n4 <= '1';
   U3 : INV_X1 port map( A => n13, ZN => n2);
   U4 : INV_X1 port map( A => n11, ZN => n3);
   U5 : OR4_X1 port map( A1 => n5, A2 => n2, A3 => n3, A4 => n114, ZN => n10);
   U6 : INV_X1 port map( A => n10, ZN => n1);
   U7 : NOR3_X4 port map( A1 => n115, A2 => SEL(1), A3 => n117, ZN => n15);
   U8 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(1), A3 => n115, ZN => n17);
   U9 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(2), A3 => n116, ZN => n14);
   U10 : NOR3_X4 port map( A1 => n117, A2 => n115, A3 => n116, ZN => n16);
   U11 : OR3_X1 port map( A1 => n117, A2 => SEL(2), A3 => n116, ZN => n13);
   U12 : OR3_X1 port map( A1 => n115, A2 => SEL(0), A3 => n116, ZN => n11);
   U13 : OR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n117, ZN => n12);
   U14 : INV_X2 port map( A => n12, ZN => n5);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => N195)
                           ;
   U16 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(150), B2 =>
                           n3, ZN => n9);
   U17 : AOI22_X1 port map( A1 => inputs(25), A2 => n5, B1 => inputs(75), B2 =>
                           n2, ZN => n8);
   U18 : AOI22_X1 port map( A1 => inputs(50), A2 => n14, B1 => inputs(125), B2 
                           => n15, ZN => n7);
   U19 : AOI22_X1 port map( A1 => inputs(175), A2 => n16, B1 => inputs(100), B2
                           => n17, ZN => n6);
   U20 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           N194);
   U21 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(151), B2 =>
                           n3, ZN => n21);
   U22 : AOI22_X1 port map( A1 => inputs(26), A2 => n5, B1 => inputs(76), B2 =>
                           n2, ZN => n20);
   U23 : AOI22_X1 port map( A1 => inputs(51), A2 => n14, B1 => inputs(126), B2 
                           => n15, ZN => n19);
   U24 : AOI22_X1 port map( A1 => inputs(176), A2 => n16, B1 => inputs(101), B2
                           => n17, ZN => n18);
   U25 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           N193);
   U26 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(152), B2 =>
                           n3, ZN => n25);
   U27 : AOI22_X1 port map( A1 => inputs(27), A2 => n5, B1 => inputs(77), B2 =>
                           n2, ZN => n24);
   U28 : AOI22_X1 port map( A1 => inputs(52), A2 => n14, B1 => inputs(127), B2 
                           => n15, ZN => n23);
   U29 : AOI22_X1 port map( A1 => inputs(177), A2 => n16, B1 => inputs(102), B2
                           => n17, ZN => n22);
   U30 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n28, A4 => n29, ZN => 
                           N192);
   U31 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(153), B2 =>
                           n3, ZN => n29);
   U32 : AOI22_X1 port map( A1 => inputs(28), A2 => n5, B1 => inputs(78), B2 =>
                           n2, ZN => n28);
   U33 : AOI22_X1 port map( A1 => inputs(53), A2 => n14, B1 => inputs(128), B2 
                           => n15, ZN => n27);
   U34 : AOI22_X1 port map( A1 => inputs(178), A2 => n16, B1 => inputs(103), B2
                           => n17, ZN => n26);
   U35 : NAND4_X1 port map( A1 => n30, A2 => n31, A3 => n32, A4 => n33, ZN => 
                           N191);
   U36 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(154), B2 =>
                           n3, ZN => n33);
   U37 : AOI22_X1 port map( A1 => inputs(29), A2 => n5, B1 => inputs(79), B2 =>
                           n2, ZN => n32);
   U38 : AOI22_X1 port map( A1 => inputs(54), A2 => n14, B1 => inputs(129), B2 
                           => n15, ZN => n31);
   U39 : AOI22_X1 port map( A1 => inputs(179), A2 => n16, B1 => inputs(104), B2
                           => n17, ZN => n30);
   U40 : NAND4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           N190);
   U41 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(155), B2 =>
                           n3, ZN => n37);
   U42 : AOI22_X1 port map( A1 => inputs(30), A2 => n5, B1 => inputs(80), B2 =>
                           n2, ZN => n36);
   U43 : AOI22_X1 port map( A1 => inputs(55), A2 => n14, B1 => inputs(130), B2 
                           => n15, ZN => n35);
   U44 : AOI22_X1 port map( A1 => inputs(180), A2 => n16, B1 => inputs(105), B2
                           => n17, ZN => n34);
   U45 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           N189);
   U46 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(156), B2 =>
                           n3, ZN => n41);
   U47 : AOI22_X1 port map( A1 => inputs(31), A2 => n5, B1 => inputs(81), B2 =>
                           n2, ZN => n40);
   U48 : AOI22_X1 port map( A1 => inputs(56), A2 => n14, B1 => inputs(131), B2 
                           => n15, ZN => n39);
   U49 : AOI22_X1 port map( A1 => inputs(181), A2 => n16, B1 => inputs(106), B2
                           => n17, ZN => n38);
   U50 : NAND4_X1 port map( A1 => n42, A2 => n43, A3 => n44, A4 => n45, ZN => 
                           N188);
   U51 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(157), B2 =>
                           n3, ZN => n45);
   U52 : AOI22_X1 port map( A1 => inputs(32), A2 => n5, B1 => inputs(82), B2 =>
                           n2, ZN => n44);
   U53 : AOI22_X1 port map( A1 => inputs(57), A2 => n14, B1 => inputs(132), B2 
                           => n15, ZN => n43);
   U54 : AOI22_X1 port map( A1 => inputs(182), A2 => n16, B1 => inputs(107), B2
                           => n17, ZN => n42);
   U55 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           N187);
   U56 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(158), B2 =>
                           n3, ZN => n49);
   U57 : AOI22_X1 port map( A1 => inputs(33), A2 => n5, B1 => inputs(83), B2 =>
                           n2, ZN => n48);
   U58 : AOI22_X1 port map( A1 => inputs(58), A2 => n14, B1 => inputs(133), B2 
                           => n15, ZN => n47);
   U59 : AOI22_X1 port map( A1 => inputs(183), A2 => n16, B1 => inputs(108), B2
                           => n17, ZN => n46);
   U60 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           N186);
   U61 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(159), B2 =>
                           n3, ZN => n53);
   U62 : AOI22_X1 port map( A1 => inputs(34), A2 => n5, B1 => inputs(84), B2 =>
                           n2, ZN => n52);
   U63 : AOI22_X1 port map( A1 => inputs(59), A2 => n14, B1 => inputs(134), B2 
                           => n15, ZN => n51);
   U64 : AOI22_X1 port map( A1 => inputs(184), A2 => n16, B1 => inputs(109), B2
                           => n17, ZN => n50);
   U65 : NAND4_X1 port map( A1 => n54, A2 => n55, A3 => n56, A4 => n57, ZN => 
                           N185);
   U66 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(160), B2 
                           => n3, ZN => n57);
   U67 : AOI22_X1 port map( A1 => inputs(35), A2 => n5, B1 => inputs(85), B2 =>
                           n2, ZN => n56);
   U68 : AOI22_X1 port map( A1 => inputs(60), A2 => n14, B1 => inputs(135), B2 
                           => n15, ZN => n55);
   U69 : AOI22_X1 port map( A1 => inputs(185), A2 => n16, B1 => inputs(110), B2
                           => n17, ZN => n54);
   U70 : NAND4_X1 port map( A1 => n58, A2 => n59, A3 => n60, A4 => n61, ZN => 
                           N184);
   U71 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(161), B2 
                           => n3, ZN => n61);
   U72 : AOI22_X1 port map( A1 => inputs(36), A2 => n5, B1 => inputs(86), B2 =>
                           n2, ZN => n60);
   U73 : AOI22_X1 port map( A1 => inputs(61), A2 => n14, B1 => inputs(136), B2 
                           => n15, ZN => n59);
   U74 : AOI22_X1 port map( A1 => inputs(186), A2 => n16, B1 => inputs(111), B2
                           => n17, ZN => n58);
   U75 : NAND4_X1 port map( A1 => n62, A2 => n63, A3 => n64, A4 => n65, ZN => 
                           N183);
   U76 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(162), B2 
                           => n3, ZN => n65);
   U77 : AOI22_X1 port map( A1 => inputs(37), A2 => n5, B1 => inputs(87), B2 =>
                           n2, ZN => n64);
   U78 : AOI22_X1 port map( A1 => inputs(62), A2 => n14, B1 => inputs(137), B2 
                           => n15, ZN => n63);
   U79 : AOI22_X1 port map( A1 => inputs(187), A2 => n16, B1 => inputs(112), B2
                           => n17, ZN => n62);
   U80 : NAND4_X1 port map( A1 => n66, A2 => n67, A3 => n68, A4 => n69, ZN => 
                           N182);
   U81 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(163), B2 
                           => n3, ZN => n69);
   U82 : AOI22_X1 port map( A1 => inputs(38), A2 => n5, B1 => inputs(88), B2 =>
                           n2, ZN => n68);
   U83 : AOI22_X1 port map( A1 => inputs(63), A2 => n14, B1 => inputs(138), B2 
                           => n15, ZN => n67);
   U84 : AOI22_X1 port map( A1 => inputs(188), A2 => n16, B1 => inputs(113), B2
                           => n17, ZN => n66);
   U85 : NAND4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           N181);
   U86 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(164), B2 
                           => n3, ZN => n73);
   U87 : AOI22_X1 port map( A1 => inputs(39), A2 => n5, B1 => inputs(89), B2 =>
                           n2, ZN => n72);
   U88 : AOI22_X1 port map( A1 => inputs(64), A2 => n14, B1 => inputs(139), B2 
                           => n15, ZN => n71);
   U89 : AOI22_X1 port map( A1 => inputs(189), A2 => n16, B1 => inputs(114), B2
                           => n17, ZN => n70);
   U90 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           N180);
   U91 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(165), B2 
                           => n3, ZN => n77);
   U92 : AOI22_X1 port map( A1 => inputs(40), A2 => n5, B1 => inputs(90), B2 =>
                           n2, ZN => n76);
   U93 : AOI22_X1 port map( A1 => inputs(65), A2 => n14, B1 => inputs(140), B2 
                           => n15, ZN => n75);
   U94 : AOI22_X1 port map( A1 => inputs(190), A2 => n16, B1 => inputs(115), B2
                           => n17, ZN => n74);
   U95 : NAND4_X1 port map( A1 => n78, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           N179);
   U96 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(166), B2 
                           => n3, ZN => n81);
   U97 : AOI22_X1 port map( A1 => inputs(41), A2 => n5, B1 => inputs(91), B2 =>
                           n2, ZN => n80);
   U98 : AOI22_X1 port map( A1 => inputs(66), A2 => n14, B1 => inputs(141), B2 
                           => n15, ZN => n79);
   U99 : AOI22_X1 port map( A1 => inputs(191), A2 => n16, B1 => inputs(116), B2
                           => n17, ZN => n78);
   U100 : NAND4_X1 port map( A1 => n82, A2 => n83, A3 => n84, A4 => n85, ZN => 
                           N178);
   U101 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(167), B2 
                           => n3, ZN => n85);
   U102 : AOI22_X1 port map( A1 => inputs(42), A2 => n5, B1 => inputs(92), B2 
                           => n2, ZN => n84);
   U103 : AOI22_X1 port map( A1 => inputs(67), A2 => n14, B1 => inputs(142), B2
                           => n15, ZN => n83);
   U104 : AOI22_X1 port map( A1 => inputs(192), A2 => n16, B1 => inputs(117), 
                           B2 => n17, ZN => n82);
   U105 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           N177);
   U106 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(168), B2 
                           => n3, ZN => n89);
   U107 : AOI22_X1 port map( A1 => inputs(43), A2 => n5, B1 => inputs(93), B2 
                           => n2, ZN => n88);
   U108 : AOI22_X1 port map( A1 => inputs(68), A2 => n14, B1 => inputs(143), B2
                           => n15, ZN => n87);
   U109 : AOI22_X1 port map( A1 => inputs(193), A2 => n16, B1 => inputs(118), 
                           B2 => n17, ZN => n86);
   U110 : NAND4_X1 port map( A1 => n90, A2 => n91, A3 => n92, A4 => n93, ZN => 
                           N176);
   U111 : AOI22_X1 port map( A1 => inputs(19), A2 => n1, B1 => inputs(169), B2 
                           => n3, ZN => n93);
   U112 : AOI22_X1 port map( A1 => inputs(44), A2 => n5, B1 => inputs(94), B2 
                           => n2, ZN => n92);
   U113 : AOI22_X1 port map( A1 => inputs(69), A2 => n14, B1 => inputs(144), B2
                           => n15, ZN => n91);
   U114 : AOI22_X1 port map( A1 => inputs(194), A2 => n16, B1 => inputs(119), 
                           B2 => n17, ZN => n90);
   U115 : NAND4_X1 port map( A1 => n94, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           N175);
   U116 : AOI22_X1 port map( A1 => inputs(20), A2 => n1, B1 => inputs(170), B2 
                           => n3, ZN => n97);
   U117 : AOI22_X1 port map( A1 => inputs(45), A2 => n5, B1 => inputs(95), B2 
                           => n2, ZN => n96);
   U118 : AOI22_X1 port map( A1 => inputs(70), A2 => n14, B1 => inputs(145), B2
                           => n15, ZN => n95);
   U119 : AOI22_X1 port map( A1 => inputs(195), A2 => n16, B1 => inputs(120), 
                           B2 => n17, ZN => n94);
   U120 : NAND4_X1 port map( A1 => n98, A2 => n99, A3 => n100, A4 => n101, ZN 
                           => N174);
   U121 : AOI22_X1 port map( A1 => inputs(21), A2 => n1, B1 => inputs(171), B2 
                           => n3, ZN => n101);
   U122 : AOI22_X1 port map( A1 => inputs(46), A2 => n5, B1 => inputs(96), B2 
                           => n2, ZN => n100);
   U123 : AOI22_X1 port map( A1 => inputs(71), A2 => n14, B1 => inputs(146), B2
                           => n15, ZN => n99);
   U124 : AOI22_X1 port map( A1 => inputs(196), A2 => n16, B1 => inputs(121), 
                           B2 => n17, ZN => n98);
   U125 : NAND4_X1 port map( A1 => n102, A2 => n103, A3 => n104, A4 => n105, ZN
                           => N173);
   U126 : AOI22_X1 port map( A1 => inputs(22), A2 => n1, B1 => inputs(172), B2 
                           => n3, ZN => n105);
   U127 : AOI22_X1 port map( A1 => inputs(47), A2 => n5, B1 => inputs(97), B2 
                           => n2, ZN => n104);
   U128 : AOI22_X1 port map( A1 => inputs(72), A2 => n14, B1 => inputs(147), B2
                           => n15, ZN => n103);
   U129 : AOI22_X1 port map( A1 => inputs(197), A2 => n16, B1 => inputs(122), 
                           B2 => n17, ZN => n102);
   U130 : NAND4_X1 port map( A1 => n106, A2 => n107, A3 => n108, A4 => n109, ZN
                           => N172);
   U131 : AOI22_X1 port map( A1 => inputs(23), A2 => n1, B1 => inputs(173), B2 
                           => n3, ZN => n109);
   U132 : AOI22_X1 port map( A1 => inputs(48), A2 => n5, B1 => inputs(98), B2 
                           => n2, ZN => n108);
   U133 : AOI22_X1 port map( A1 => inputs(73), A2 => n14, B1 => inputs(148), B2
                           => n15, ZN => n107);
   U134 : AOI22_X1 port map( A1 => inputs(198), A2 => n16, B1 => inputs(123), 
                           B2 => n17, ZN => n106);
   U135 : NAND4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN
                           => N171);
   U136 : AOI22_X1 port map( A1 => inputs(24), A2 => n1, B1 => inputs(174), B2 
                           => n3, ZN => n113);
   U137 : OR4_X1 port map( A1 => n17, A2 => n16, A3 => n15, A4 => n14, ZN => 
                           n114);
   U138 : AOI22_X1 port map( A1 => inputs(49), A2 => n5, B1 => inputs(99), B2 
                           => n2, ZN => n112);
   U139 : AOI22_X1 port map( A1 => inputs(74), A2 => n14, B1 => inputs(149), B2
                           => n15, ZN => n111);
   U141 : AOI22_X1 port map( A1 => inputs(199), A2 => n16, B1 => inputs(124), 
                           B2 => n17, ZN => n110);
   U142 : INV_X1 port map( A => SEL(1), ZN => n116);
   U143 : INV_X1 port map( A => SEL(2), ZN => n115);
   U144 : INV_X1 port map( A => SEL(0), ZN => n117);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT23 is

   port( a, b : in std_logic_vector (22 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (23 downto 0));

end adder_NBIT23;

architecture SYN_beh of adder_NBIT23 is

   component adder_NBIT23_DW01_add_0
      port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (23 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3353 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT23_DW01_add_0 port map( A(23) => a(22), 
                           A(22) => a(22), A(21) => a(21), A(20) => a(20), 
                           A(19) => a(19), A(18) => a(18), A(17) => a(17), 
                           A(16) => a(16), A(15) => a(15), A(14) => a(14), 
                           A(13) => a(13), A(12) => a(12), A(11) => a(11), 
                           A(10) => a(10), A(9) => a(9), A(8) => a(8), A(7) => 
                           a(7), A(6) => a(6), A(5) => a(5), A(4) => a(4), A(3)
                           => a(3), A(2) => a(2), A(1) => a(1), A(0) => a(0), 
                           B(23) => b(22), B(22) => b(22), B(21) => b(21), 
                           B(20) => b(20), B(19) => b(19), B(18) => b(18), 
                           B(17) => b(17), B(16) => b(16), B(15) => b(15), 
                           B(14) => b(14), B(13) => b(13), B(12) => b(12), 
                           B(11) => b(11), B(10) => b(10), B(9) => b(9), B(8) 
                           => b(8), B(7) => b(7), B(6) => b(6), B(5) => b(5), 
                           B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1) => 
                           b(1), B(0) => b(0), CI => cin, SUM(23) => s(23), 
                           SUM(22) => s(22), SUM(21) => s(21), SUM(20) => s(20)
                           , SUM(19) => s(19), SUM(18) => s(18), SUM(17) => 
                           s(17), SUM(16) => s(16), SUM(15) => s(15), SUM(14) 
                           => s(14), SUM(13) => s(13), SUM(12) => s(12), 
                           SUM(11) => s(11), SUM(10) => s(10), SUM(9) => s(9), 
                           SUM(8) => s(8), SUM(7) => s(7), SUM(6) => s(6), 
                           SUM(5) => s(5), SUM(4) => s(4), SUM(3) => s(3), 
                           SUM(2) => s(2), SUM(1) => s(1), SUM(0) => s(0), CO 
                           => n_3353);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N23_Z3 is

   port( inputs : in std_logic_vector (0 to 183);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (22 downto 0));

end MUX_zbit_nbit_N23_Z3;

architecture SYN_beh of MUX_zbit_nbit_N23_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, 
      N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, 
      n4, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106 : std_logic;

begin
   
   Y_reg_22_inst : DLH_X1 port map( G => n4, D => N181, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n4, D => N180, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N179, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N178, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N177, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N176, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N175, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N174, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N173, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N172, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N171, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N170, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N169, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N168, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N167, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N166, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N165, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N164, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N163, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N162, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N161, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N160, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N159, Q => Y(0));
   n4 <= '1';
   U3 : OR4_X1 port map( A1 => n9, A2 => n10, A3 => n8, A4 => n103, ZN => n7);
   U4 : INV_X1 port map( A => n7, ZN => n1);
   U5 : NOR3_X4 port map( A1 => n104, A2 => SEL(1), A3 => n106, ZN => n12);
   U6 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(1), A3 => n104, ZN => n14);
   U7 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(2), A3 => n105, ZN => n11);
   U8 : NOR3_X4 port map( A1 => n106, A2 => n104, A3 => n105, ZN => n13);
   U9 : NOR3_X4 port map( A1 => n106, A2 => SEL(2), A3 => n105, ZN => n10);
   U10 : NOR3_X4 port map( A1 => n104, A2 => SEL(0), A3 => n105, ZN => n8);
   U11 : NOR3_X4 port map( A1 => SEL(1), A2 => SEL(2), A3 => n106, ZN => n9);
   U12 : NAND4_X1 port map( A1 => n2, A2 => n3, A3 => n5, A4 => n6, ZN => N181)
                           ;
   U13 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(138), B2 =>
                           n8, ZN => n6);
   U14 : AOI22_X1 port map( A1 => inputs(23), A2 => n9, B1 => inputs(69), B2 =>
                           n10, ZN => n5);
   U15 : AOI22_X1 port map( A1 => inputs(46), A2 => n11, B1 => inputs(115), B2 
                           => n12, ZN => n3);
   U16 : AOI22_X1 port map( A1 => inputs(161), A2 => n13, B1 => inputs(92), B2 
                           => n14, ZN => n2);
   U17 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           N180);
   U18 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(139), B2 =>
                           n8, ZN => n18);
   U19 : AOI22_X1 port map( A1 => inputs(24), A2 => n9, B1 => inputs(70), B2 =>
                           n10, ZN => n17);
   U20 : AOI22_X1 port map( A1 => inputs(47), A2 => n11, B1 => inputs(116), B2 
                           => n12, ZN => n16);
   U21 : AOI22_X1 port map( A1 => inputs(162), A2 => n13, B1 => inputs(93), B2 
                           => n14, ZN => n15);
   U22 : NAND4_X1 port map( A1 => n19, A2 => n20, A3 => n21, A4 => n22, ZN => 
                           N179);
   U23 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(140), B2 =>
                           n8, ZN => n22);
   U24 : AOI22_X1 port map( A1 => inputs(25), A2 => n9, B1 => inputs(71), B2 =>
                           n10, ZN => n21);
   U25 : AOI22_X1 port map( A1 => inputs(48), A2 => n11, B1 => inputs(117), B2 
                           => n12, ZN => n20);
   U26 : AOI22_X1 port map( A1 => inputs(163), A2 => n13, B1 => inputs(94), B2 
                           => n14, ZN => n19);
   U27 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           N178);
   U28 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(141), B2 =>
                           n8, ZN => n26);
   U29 : AOI22_X1 port map( A1 => inputs(26), A2 => n9, B1 => inputs(72), B2 =>
                           n10, ZN => n25);
   U30 : AOI22_X1 port map( A1 => inputs(49), A2 => n11, B1 => inputs(118), B2 
                           => n12, ZN => n24);
   U31 : AOI22_X1 port map( A1 => inputs(164), A2 => n13, B1 => inputs(95), B2 
                           => n14, ZN => n23);
   U32 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n30, ZN => 
                           N177);
   U33 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(142), B2 =>
                           n8, ZN => n30);
   U34 : AOI22_X1 port map( A1 => inputs(27), A2 => n9, B1 => inputs(73), B2 =>
                           n10, ZN => n29);
   U35 : AOI22_X1 port map( A1 => inputs(50), A2 => n11, B1 => inputs(119), B2 
                           => n12, ZN => n28);
   U36 : AOI22_X1 port map( A1 => inputs(165), A2 => n13, B1 => inputs(96), B2 
                           => n14, ZN => n27);
   U37 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           N176);
   U38 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(143), B2 =>
                           n8, ZN => n34);
   U39 : AOI22_X1 port map( A1 => inputs(28), A2 => n9, B1 => inputs(74), B2 =>
                           n10, ZN => n33);
   U40 : AOI22_X1 port map( A1 => inputs(51), A2 => n11, B1 => inputs(120), B2 
                           => n12, ZN => n32);
   U41 : AOI22_X1 port map( A1 => inputs(166), A2 => n13, B1 => inputs(97), B2 
                           => n14, ZN => n31);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           N175);
   U43 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(144), B2 =>
                           n8, ZN => n38);
   U44 : AOI22_X1 port map( A1 => inputs(29), A2 => n9, B1 => inputs(75), B2 =>
                           n10, ZN => n37);
   U45 : AOI22_X1 port map( A1 => inputs(52), A2 => n11, B1 => inputs(121), B2 
                           => n12, ZN => n36);
   U46 : AOI22_X1 port map( A1 => inputs(167), A2 => n13, B1 => inputs(98), B2 
                           => n14, ZN => n35);
   U47 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           N174);
   U48 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(145), B2 =>
                           n8, ZN => n42);
   U49 : AOI22_X1 port map( A1 => inputs(30), A2 => n9, B1 => inputs(76), B2 =>
                           n10, ZN => n41);
   U50 : AOI22_X1 port map( A1 => inputs(53), A2 => n11, B1 => inputs(122), B2 
                           => n12, ZN => n40);
   U51 : AOI22_X1 port map( A1 => inputs(168), A2 => n13, B1 => inputs(99), B2 
                           => n14, ZN => n39);
   U52 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           N173);
   U53 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(146), B2 =>
                           n8, ZN => n46);
   U54 : AOI22_X1 port map( A1 => inputs(31), A2 => n9, B1 => inputs(77), B2 =>
                           n10, ZN => n45);
   U55 : AOI22_X1 port map( A1 => inputs(54), A2 => n11, B1 => inputs(123), B2 
                           => n12, ZN => n44);
   U56 : AOI22_X1 port map( A1 => inputs(169), A2 => n13, B1 => inputs(100), B2
                           => n14, ZN => n43);
   U57 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           N172);
   U58 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(147), B2 =>
                           n8, ZN => n50);
   U59 : AOI22_X1 port map( A1 => inputs(32), A2 => n9, B1 => inputs(78), B2 =>
                           n10, ZN => n49);
   U60 : AOI22_X1 port map( A1 => inputs(55), A2 => n11, B1 => inputs(124), B2 
                           => n12, ZN => n48);
   U61 : AOI22_X1 port map( A1 => inputs(170), A2 => n13, B1 => inputs(101), B2
                           => n14, ZN => n47);
   U62 : NAND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           N171);
   U63 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(148), B2 
                           => n8, ZN => n54);
   U64 : AOI22_X1 port map( A1 => inputs(33), A2 => n9, B1 => inputs(79), B2 =>
                           n10, ZN => n53);
   U65 : AOI22_X1 port map( A1 => inputs(56), A2 => n11, B1 => inputs(125), B2 
                           => n12, ZN => n52);
   U66 : AOI22_X1 port map( A1 => inputs(171), A2 => n13, B1 => inputs(102), B2
                           => n14, ZN => n51);
   U67 : NAND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           N170);
   U68 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(149), B2 
                           => n8, ZN => n58);
   U69 : AOI22_X1 port map( A1 => inputs(34), A2 => n9, B1 => inputs(80), B2 =>
                           n10, ZN => n57);
   U70 : AOI22_X1 port map( A1 => inputs(57), A2 => n11, B1 => inputs(126), B2 
                           => n12, ZN => n56);
   U71 : AOI22_X1 port map( A1 => inputs(172), A2 => n13, B1 => inputs(103), B2
                           => n14, ZN => n55);
   U72 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           N169);
   U73 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(150), B2 
                           => n8, ZN => n62);
   U74 : AOI22_X1 port map( A1 => inputs(35), A2 => n9, B1 => inputs(81), B2 =>
                           n10, ZN => n61);
   U75 : AOI22_X1 port map( A1 => inputs(58), A2 => n11, B1 => inputs(127), B2 
                           => n12, ZN => n60);
   U76 : AOI22_X1 port map( A1 => inputs(173), A2 => n13, B1 => inputs(104), B2
                           => n14, ZN => n59);
   U77 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           N168);
   U78 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(151), B2 
                           => n8, ZN => n66);
   U79 : AOI22_X1 port map( A1 => inputs(36), A2 => n9, B1 => inputs(82), B2 =>
                           n10, ZN => n65);
   U80 : AOI22_X1 port map( A1 => inputs(59), A2 => n11, B1 => inputs(128), B2 
                           => n12, ZN => n64);
   U81 : AOI22_X1 port map( A1 => inputs(174), A2 => n13, B1 => inputs(105), B2
                           => n14, ZN => n63);
   U82 : NAND4_X1 port map( A1 => n67, A2 => n68, A3 => n69, A4 => n70, ZN => 
                           N167);
   U83 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(152), B2 
                           => n8, ZN => n70);
   U84 : AOI22_X1 port map( A1 => inputs(37), A2 => n9, B1 => inputs(83), B2 =>
                           n10, ZN => n69);
   U85 : AOI22_X1 port map( A1 => inputs(60), A2 => n11, B1 => inputs(129), B2 
                           => n12, ZN => n68);
   U86 : AOI22_X1 port map( A1 => inputs(175), A2 => n13, B1 => inputs(106), B2
                           => n14, ZN => n67);
   U87 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           N166);
   U88 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(153), B2 
                           => n8, ZN => n74);
   U89 : AOI22_X1 port map( A1 => inputs(38), A2 => n9, B1 => inputs(84), B2 =>
                           n10, ZN => n73);
   U90 : AOI22_X1 port map( A1 => inputs(61), A2 => n11, B1 => inputs(130), B2 
                           => n12, ZN => n72);
   U91 : AOI22_X1 port map( A1 => inputs(176), A2 => n13, B1 => inputs(107), B2
                           => n14, ZN => n71);
   U92 : NAND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           N165);
   U93 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(154), B2 
                           => n8, ZN => n78);
   U94 : AOI22_X1 port map( A1 => inputs(39), A2 => n9, B1 => inputs(85), B2 =>
                           n10, ZN => n77);
   U95 : AOI22_X1 port map( A1 => inputs(62), A2 => n11, B1 => inputs(131), B2 
                           => n12, ZN => n76);
   U96 : AOI22_X1 port map( A1 => inputs(177), A2 => n13, B1 => inputs(108), B2
                           => n14, ZN => n75);
   U97 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           N164);
   U98 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(155), B2 
                           => n8, ZN => n82);
   U99 : AOI22_X1 port map( A1 => inputs(40), A2 => n9, B1 => inputs(86), B2 =>
                           n10, ZN => n81);
   U100 : AOI22_X1 port map( A1 => inputs(63), A2 => n11, B1 => inputs(132), B2
                           => n12, ZN => n80);
   U101 : AOI22_X1 port map( A1 => inputs(178), A2 => n13, B1 => inputs(109), 
                           B2 => n14, ZN => n79);
   U102 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           N163);
   U103 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(156), B2 
                           => n8, ZN => n86);
   U104 : AOI22_X1 port map( A1 => inputs(41), A2 => n9, B1 => inputs(87), B2 
                           => n10, ZN => n85);
   U105 : AOI22_X1 port map( A1 => inputs(64), A2 => n11, B1 => inputs(133), B2
                           => n12, ZN => n84);
   U106 : AOI22_X1 port map( A1 => inputs(179), A2 => n13, B1 => inputs(110), 
                           B2 => n14, ZN => n83);
   U107 : NAND4_X1 port map( A1 => n87, A2 => n88, A3 => n89, A4 => n90, ZN => 
                           N162);
   U108 : AOI22_X1 port map( A1 => inputs(19), A2 => n1, B1 => inputs(157), B2 
                           => n8, ZN => n90);
   U109 : AOI22_X1 port map( A1 => inputs(42), A2 => n9, B1 => inputs(88), B2 
                           => n10, ZN => n89);
   U110 : AOI22_X1 port map( A1 => inputs(65), A2 => n11, B1 => inputs(134), B2
                           => n12, ZN => n88);
   U111 : AOI22_X1 port map( A1 => inputs(180), A2 => n13, B1 => inputs(111), 
                           B2 => n14, ZN => n87);
   U112 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           N161);
   U113 : AOI22_X1 port map( A1 => inputs(20), A2 => n1, B1 => inputs(158), B2 
                           => n8, ZN => n94);
   U114 : AOI22_X1 port map( A1 => inputs(43), A2 => n9, B1 => inputs(89), B2 
                           => n10, ZN => n93);
   U115 : AOI22_X1 port map( A1 => inputs(66), A2 => n11, B1 => inputs(135), B2
                           => n12, ZN => n92);
   U116 : AOI22_X1 port map( A1 => inputs(181), A2 => n13, B1 => inputs(112), 
                           B2 => n14, ZN => n91);
   U117 : NAND4_X1 port map( A1 => n95, A2 => n96, A3 => n97, A4 => n98, ZN => 
                           N160);
   U118 : AOI22_X1 port map( A1 => inputs(21), A2 => n1, B1 => inputs(159), B2 
                           => n8, ZN => n98);
   U119 : AOI22_X1 port map( A1 => inputs(44), A2 => n9, B1 => inputs(90), B2 
                           => n10, ZN => n97);
   U120 : AOI22_X1 port map( A1 => inputs(67), A2 => n11, B1 => inputs(136), B2
                           => n12, ZN => n96);
   U121 : AOI22_X1 port map( A1 => inputs(182), A2 => n13, B1 => inputs(113), 
                           B2 => n14, ZN => n95);
   U122 : NAND4_X1 port map( A1 => n99, A2 => n100, A3 => n101, A4 => n102, ZN 
                           => N159);
   U123 : AOI22_X1 port map( A1 => inputs(22), A2 => n1, B1 => inputs(160), B2 
                           => n8, ZN => n102);
   U124 : OR4_X1 port map( A1 => n14, A2 => n13, A3 => n12, A4 => n11, ZN => 
                           n103);
   U125 : AOI22_X1 port map( A1 => inputs(45), A2 => n9, B1 => inputs(91), B2 
                           => n10, ZN => n101);
   U126 : AOI22_X1 port map( A1 => inputs(68), A2 => n11, B1 => inputs(137), B2
                           => n12, ZN => n100);
   U127 : AOI22_X1 port map( A1 => inputs(183), A2 => n13, B1 => inputs(114), 
                           B2 => n14, ZN => n99);
   U128 : INV_X1 port map( A => SEL(1), ZN => n105);
   U129 : INV_X1 port map( A => SEL(2), ZN => n104);
   U131 : INV_X1 port map( A => SEL(0), ZN => n106);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT21 is

   port( a, b : in std_logic_vector (20 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (21 downto 0));

end adder_NBIT21;

architecture SYN_beh of adder_NBIT21 is

   component adder_NBIT21_DW01_add_0
      port( A, B : in std_logic_vector (21 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (21 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3354 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT21_DW01_add_0 port map( A(21) => a(20), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), B(21) => b(20), B(20) => b(20), 
                           B(19) => b(19), B(18) => b(18), B(17) => b(17), 
                           B(16) => b(16), B(15) => b(15), B(14) => b(14), 
                           B(13) => b(13), B(12) => b(12), B(11) => b(11), 
                           B(10) => b(10), B(9) => b(9), B(8) => b(8), B(7) => 
                           b(7), B(6) => b(6), B(5) => b(5), B(4) => b(4), B(3)
                           => b(3), B(2) => b(2), B(1) => b(1), B(0) => b(0), 
                           CI => cin, SUM(21) => s(21), SUM(20) => s(20), 
                           SUM(19) => s(19), SUM(18) => s(18), SUM(17) => s(17)
                           , SUM(16) => s(16), SUM(15) => s(15), SUM(14) => 
                           s(14), SUM(13) => s(13), SUM(12) => s(12), SUM(11) 
                           => s(11), SUM(10) => s(10), SUM(9) => s(9), SUM(8) 
                           => s(8), SUM(7) => s(7), SUM(6) => s(6), SUM(5) => 
                           s(5), SUM(4) => s(4), SUM(3) => s(3), SUM(2) => s(2)
                           , SUM(1) => s(1), SUM(0) => s(0), CO => n_3354);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N21_Z3 is

   port( inputs : in std_logic_vector (0 to 167);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (20 downto 0));

end MUX_zbit_nbit_N21_Z3;

architecture SYN_beh of MUX_zbit_nbit_N21_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, 
      N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, n4, n1, n2, 
      n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98 : std_logic;

begin
   
   Y_reg_20_inst : DLH_X1 port map( G => n4, D => N167, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n4, D => N166, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N165, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N164, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N163, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N162, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N161, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N160, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N159, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N158, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N157, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N156, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N155, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N154, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N153, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N152, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N151, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N150, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N149, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N148, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N147, Q => Y(0));
   n4 <= '1';
   U3 : OR4_X1 port map( A1 => n9, A2 => n10, A3 => n8, A4 => n95, ZN => n7);
   U4 : INV_X1 port map( A => n7, ZN => n1);
   U5 : NOR3_X4 port map( A1 => n96, A2 => SEL(1), A3 => n98, ZN => n12);
   U6 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(1), A3 => n96, ZN => n14);
   U7 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(2), A3 => n97, ZN => n11);
   U8 : NOR3_X4 port map( A1 => n98, A2 => n96, A3 => n97, ZN => n13);
   U9 : NOR3_X4 port map( A1 => n98, A2 => SEL(2), A3 => n97, ZN => n10);
   U10 : NOR3_X4 port map( A1 => n96, A2 => SEL(0), A3 => n97, ZN => n8);
   U11 : NOR3_X4 port map( A1 => SEL(1), A2 => SEL(2), A3 => n98, ZN => n9);
   U12 : NAND4_X1 port map( A1 => n2, A2 => n3, A3 => n5, A4 => n6, ZN => N167)
                           ;
   U13 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(126), B2 =>
                           n8, ZN => n6);
   U14 : AOI22_X1 port map( A1 => inputs(21), A2 => n9, B1 => inputs(63), B2 =>
                           n10, ZN => n5);
   U15 : AOI22_X1 port map( A1 => inputs(42), A2 => n11, B1 => inputs(105), B2 
                           => n12, ZN => n3);
   U16 : AOI22_X1 port map( A1 => inputs(147), A2 => n13, B1 => inputs(84), B2 
                           => n14, ZN => n2);
   U17 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           N166);
   U18 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(127), B2 =>
                           n8, ZN => n18);
   U19 : AOI22_X1 port map( A1 => inputs(22), A2 => n9, B1 => inputs(64), B2 =>
                           n10, ZN => n17);
   U20 : AOI22_X1 port map( A1 => inputs(43), A2 => n11, B1 => inputs(106), B2 
                           => n12, ZN => n16);
   U21 : AOI22_X1 port map( A1 => inputs(148), A2 => n13, B1 => inputs(85), B2 
                           => n14, ZN => n15);
   U22 : NAND4_X1 port map( A1 => n19, A2 => n20, A3 => n21, A4 => n22, ZN => 
                           N165);
   U23 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(128), B2 =>
                           n8, ZN => n22);
   U24 : AOI22_X1 port map( A1 => inputs(23), A2 => n9, B1 => inputs(65), B2 =>
                           n10, ZN => n21);
   U25 : AOI22_X1 port map( A1 => inputs(44), A2 => n11, B1 => inputs(107), B2 
                           => n12, ZN => n20);
   U26 : AOI22_X1 port map( A1 => inputs(149), A2 => n13, B1 => inputs(86), B2 
                           => n14, ZN => n19);
   U27 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           N164);
   U28 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(129), B2 =>
                           n8, ZN => n26);
   U29 : AOI22_X1 port map( A1 => inputs(24), A2 => n9, B1 => inputs(66), B2 =>
                           n10, ZN => n25);
   U30 : AOI22_X1 port map( A1 => inputs(45), A2 => n11, B1 => inputs(108), B2 
                           => n12, ZN => n24);
   U31 : AOI22_X1 port map( A1 => inputs(150), A2 => n13, B1 => inputs(87), B2 
                           => n14, ZN => n23);
   U32 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n30, ZN => 
                           N163);
   U33 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(130), B2 =>
                           n8, ZN => n30);
   U34 : AOI22_X1 port map( A1 => inputs(25), A2 => n9, B1 => inputs(67), B2 =>
                           n10, ZN => n29);
   U35 : AOI22_X1 port map( A1 => inputs(46), A2 => n11, B1 => inputs(109), B2 
                           => n12, ZN => n28);
   U36 : AOI22_X1 port map( A1 => inputs(151), A2 => n13, B1 => inputs(88), B2 
                           => n14, ZN => n27);
   U37 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           N162);
   U38 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(131), B2 =>
                           n8, ZN => n34);
   U39 : AOI22_X1 port map( A1 => inputs(26), A2 => n9, B1 => inputs(68), B2 =>
                           n10, ZN => n33);
   U40 : AOI22_X1 port map( A1 => inputs(47), A2 => n11, B1 => inputs(110), B2 
                           => n12, ZN => n32);
   U41 : AOI22_X1 port map( A1 => inputs(152), A2 => n13, B1 => inputs(89), B2 
                           => n14, ZN => n31);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           N161);
   U43 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(132), B2 =>
                           n8, ZN => n38);
   U44 : AOI22_X1 port map( A1 => inputs(27), A2 => n9, B1 => inputs(69), B2 =>
                           n10, ZN => n37);
   U45 : AOI22_X1 port map( A1 => inputs(48), A2 => n11, B1 => inputs(111), B2 
                           => n12, ZN => n36);
   U46 : AOI22_X1 port map( A1 => inputs(153), A2 => n13, B1 => inputs(90), B2 
                           => n14, ZN => n35);
   U47 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           N160);
   U48 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(133), B2 =>
                           n8, ZN => n42);
   U49 : AOI22_X1 port map( A1 => inputs(28), A2 => n9, B1 => inputs(70), B2 =>
                           n10, ZN => n41);
   U50 : AOI22_X1 port map( A1 => inputs(49), A2 => n11, B1 => inputs(112), B2 
                           => n12, ZN => n40);
   U51 : AOI22_X1 port map( A1 => inputs(154), A2 => n13, B1 => inputs(91), B2 
                           => n14, ZN => n39);
   U52 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           N159);
   U53 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(134), B2 =>
                           n8, ZN => n46);
   U54 : AOI22_X1 port map( A1 => inputs(29), A2 => n9, B1 => inputs(71), B2 =>
                           n10, ZN => n45);
   U55 : AOI22_X1 port map( A1 => inputs(50), A2 => n11, B1 => inputs(113), B2 
                           => n12, ZN => n44);
   U56 : AOI22_X1 port map( A1 => inputs(155), A2 => n13, B1 => inputs(92), B2 
                           => n14, ZN => n43);
   U57 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           N158);
   U58 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(135), B2 =>
                           n8, ZN => n50);
   U59 : AOI22_X1 port map( A1 => inputs(30), A2 => n9, B1 => inputs(72), B2 =>
                           n10, ZN => n49);
   U60 : AOI22_X1 port map( A1 => inputs(51), A2 => n11, B1 => inputs(114), B2 
                           => n12, ZN => n48);
   U61 : AOI22_X1 port map( A1 => inputs(156), A2 => n13, B1 => inputs(93), B2 
                           => n14, ZN => n47);
   U62 : NAND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           N157);
   U63 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(136), B2 
                           => n8, ZN => n54);
   U64 : AOI22_X1 port map( A1 => inputs(31), A2 => n9, B1 => inputs(73), B2 =>
                           n10, ZN => n53);
   U65 : AOI22_X1 port map( A1 => inputs(52), A2 => n11, B1 => inputs(115), B2 
                           => n12, ZN => n52);
   U66 : AOI22_X1 port map( A1 => inputs(157), A2 => n13, B1 => inputs(94), B2 
                           => n14, ZN => n51);
   U67 : NAND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           N156);
   U68 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(137), B2 
                           => n8, ZN => n58);
   U69 : AOI22_X1 port map( A1 => inputs(32), A2 => n9, B1 => inputs(74), B2 =>
                           n10, ZN => n57);
   U70 : AOI22_X1 port map( A1 => inputs(53), A2 => n11, B1 => inputs(116), B2 
                           => n12, ZN => n56);
   U71 : AOI22_X1 port map( A1 => inputs(158), A2 => n13, B1 => inputs(95), B2 
                           => n14, ZN => n55);
   U72 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           N155);
   U73 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(138), B2 
                           => n8, ZN => n62);
   U74 : AOI22_X1 port map( A1 => inputs(33), A2 => n9, B1 => inputs(75), B2 =>
                           n10, ZN => n61);
   U75 : AOI22_X1 port map( A1 => inputs(54), A2 => n11, B1 => inputs(117), B2 
                           => n12, ZN => n60);
   U76 : AOI22_X1 port map( A1 => inputs(159), A2 => n13, B1 => inputs(96), B2 
                           => n14, ZN => n59);
   U77 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           N154);
   U78 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(139), B2 
                           => n8, ZN => n66);
   U79 : AOI22_X1 port map( A1 => inputs(34), A2 => n9, B1 => inputs(76), B2 =>
                           n10, ZN => n65);
   U80 : AOI22_X1 port map( A1 => inputs(55), A2 => n11, B1 => inputs(118), B2 
                           => n12, ZN => n64);
   U81 : AOI22_X1 port map( A1 => inputs(160), A2 => n13, B1 => inputs(97), B2 
                           => n14, ZN => n63);
   U82 : NAND4_X1 port map( A1 => n67, A2 => n68, A3 => n69, A4 => n70, ZN => 
                           N153);
   U83 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(140), B2 
                           => n8, ZN => n70);
   U84 : AOI22_X1 port map( A1 => inputs(35), A2 => n9, B1 => inputs(77), B2 =>
                           n10, ZN => n69);
   U85 : AOI22_X1 port map( A1 => inputs(56), A2 => n11, B1 => inputs(119), B2 
                           => n12, ZN => n68);
   U86 : AOI22_X1 port map( A1 => inputs(161), A2 => n13, B1 => inputs(98), B2 
                           => n14, ZN => n67);
   U87 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           N152);
   U88 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(141), B2 
                           => n8, ZN => n74);
   U89 : AOI22_X1 port map( A1 => inputs(36), A2 => n9, B1 => inputs(78), B2 =>
                           n10, ZN => n73);
   U90 : AOI22_X1 port map( A1 => inputs(57), A2 => n11, B1 => inputs(120), B2 
                           => n12, ZN => n72);
   U91 : AOI22_X1 port map( A1 => inputs(162), A2 => n13, B1 => inputs(99), B2 
                           => n14, ZN => n71);
   U92 : NAND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           N151);
   U93 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(142), B2 
                           => n8, ZN => n78);
   U94 : AOI22_X1 port map( A1 => inputs(37), A2 => n9, B1 => inputs(79), B2 =>
                           n10, ZN => n77);
   U95 : AOI22_X1 port map( A1 => inputs(58), A2 => n11, B1 => inputs(121), B2 
                           => n12, ZN => n76);
   U96 : AOI22_X1 port map( A1 => inputs(163), A2 => n13, B1 => inputs(100), B2
                           => n14, ZN => n75);
   U97 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           N150);
   U98 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(143), B2 
                           => n8, ZN => n82);
   U99 : AOI22_X1 port map( A1 => inputs(38), A2 => n9, B1 => inputs(80), B2 =>
                           n10, ZN => n81);
   U100 : AOI22_X1 port map( A1 => inputs(59), A2 => n11, B1 => inputs(122), B2
                           => n12, ZN => n80);
   U101 : AOI22_X1 port map( A1 => inputs(164), A2 => n13, B1 => inputs(101), 
                           B2 => n14, ZN => n79);
   U102 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           N149);
   U103 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(144), B2 
                           => n8, ZN => n86);
   U104 : AOI22_X1 port map( A1 => inputs(39), A2 => n9, B1 => inputs(81), B2 
                           => n10, ZN => n85);
   U105 : AOI22_X1 port map( A1 => inputs(60), A2 => n11, B1 => inputs(123), B2
                           => n12, ZN => n84);
   U106 : AOI22_X1 port map( A1 => inputs(165), A2 => n13, B1 => inputs(102), 
                           B2 => n14, ZN => n83);
   U107 : NAND4_X1 port map( A1 => n87, A2 => n88, A3 => n89, A4 => n90, ZN => 
                           N148);
   U108 : AOI22_X1 port map( A1 => inputs(19), A2 => n1, B1 => inputs(145), B2 
                           => n8, ZN => n90);
   U109 : AOI22_X1 port map( A1 => inputs(40), A2 => n9, B1 => inputs(82), B2 
                           => n10, ZN => n89);
   U110 : AOI22_X1 port map( A1 => inputs(61), A2 => n11, B1 => inputs(124), B2
                           => n12, ZN => n88);
   U111 : AOI22_X1 port map( A1 => inputs(166), A2 => n13, B1 => inputs(103), 
                           B2 => n14, ZN => n87);
   U112 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           N147);
   U113 : AOI22_X1 port map( A1 => inputs(20), A2 => n1, B1 => inputs(146), B2 
                           => n8, ZN => n94);
   U114 : OR4_X1 port map( A1 => n14, A2 => n13, A3 => n12, A4 => n11, ZN => 
                           n95);
   U115 : AOI22_X1 port map( A1 => inputs(41), A2 => n9, B1 => inputs(83), B2 
                           => n10, ZN => n93);
   U116 : AOI22_X1 port map( A1 => inputs(62), A2 => n11, B1 => inputs(125), B2
                           => n12, ZN => n92);
   U117 : AOI22_X1 port map( A1 => inputs(167), A2 => n13, B1 => inputs(104), 
                           B2 => n14, ZN => n91);
   U118 : INV_X1 port map( A => SEL(1), ZN => n97);
   U119 : INV_X1 port map( A => SEL(2), ZN => n96);
   U121 : INV_X1 port map( A => SEL(0), ZN => n98);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n249_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);  Q
         : out std_logic_vector (248 downto 0));

end reg_nbit_n249_0;

architecture SYN_struc of reg_nbit_n249_0 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1502
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1503
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1504
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1505
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1506
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1507
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1508
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1509
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1510
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1511
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1512
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1513
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1514
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1515
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1516
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1517
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1518
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1519
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1520
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1521
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1522
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1523
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1524
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1525
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1526
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1527
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1528
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1529
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1530
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1531
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1532
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1533
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1534
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1535
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1536
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1537
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1538
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1539
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1540
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1541
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1542
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1543
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1544
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1545
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1546
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1547
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1548
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1549
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1550
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1551
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1552
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1553
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1554
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1555
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1556
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1557
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1558
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1559
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1560
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1561
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1562
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1563
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1564
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1565
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1566
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1567
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1568
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1569
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1570
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1571
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1572
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1573
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1574
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1575
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1576
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1577
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1578
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1579
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1580
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1581
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1582
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1583
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1584
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1585
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1586
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1587
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1588
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1589
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1590
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1591
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1592
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1593
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1594
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1595
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1596
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1597
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1598
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1599
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1600
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1601
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1602
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1603
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1604
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1605
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1606
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1607
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1608
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1609
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1610
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1611
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1612
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1613
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1614
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1615
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1616
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1617
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1618
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1619
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1620
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1621
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1622
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1623
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1624
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1625
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1626
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1627
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1628
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1629
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1630
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1631
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1632
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1633
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1634
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1635
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1636
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1637
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1638
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1639
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1640
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1641
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1642
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1643
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1644
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1645
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1646
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1647
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1648
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1649
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1650
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1651
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1652
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1653
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1654
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1655
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1656
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1657
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1658
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1659
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1660
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1661
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1662
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1663
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1664
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1665
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1666
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1667
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1668
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1669
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1670
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1671
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1672
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1673
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1674
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1675
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1676
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1677
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1678
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1679
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1680
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1681
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1682
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1683
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1684
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1685
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1686
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1687
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1688
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1689
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1690
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1691
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1692
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1693
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1694
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1695
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1696
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1697
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1698
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1699
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1700
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1701
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1702
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1703
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1704
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1705
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1706
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1707
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1708
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1709
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1710
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1711
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1712
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1713
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1714
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1715
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1716
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1717
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1718
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1719
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1720
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1721
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1722
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1723
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1724
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1725
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1726
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1727
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1728
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1729
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1730
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1731
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1732
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1733
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1734
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1735
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1736
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1737
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1738
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1739
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1740
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1741
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1742
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1743
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1744
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1745
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1746
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1747
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1748
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1749
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1750
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   
   D_I_0 : FD_1750 port map( D => d(0), CK => n34, RESET => n7, Q => Q(0));
   D_I_1 : FD_1749 port map( D => d(1), CK => n34, RESET => n7, Q => Q(1));
   D_I_2 : FD_1748 port map( D => d(2), CK => n34, RESET => n7, Q => Q(2));
   D_I_3 : FD_1747 port map( D => d(3), CK => n34, RESET => n7, Q => Q(3));
   D_I_4 : FD_1746 port map( D => d(4), CK => n34, RESET => n7, Q => Q(4));
   D_I_5 : FD_1745 port map( D => d(5), CK => n34, RESET => n7, Q => Q(5));
   D_I_6 : FD_1744 port map( D => d(6), CK => n34, RESET => n7, Q => Q(6));
   D_I_7 : FD_1743 port map( D => d(7), CK => n34, RESET => n7, Q => Q(7));
   D_I_8 : FD_1742 port map( D => d(8), CK => n34, RESET => n7, Q => Q(8));
   D_I_9 : FD_1741 port map( D => d(9), CK => n34, RESET => n7, Q => Q(9));
   D_I_10 : FD_1740 port map( D => d(10), CK => n34, RESET => n7, Q => Q(10));
   D_I_11 : FD_1739 port map( D => d(11), CK => n35, RESET => n7, Q => Q(11));
   D_I_12 : FD_1738 port map( D => d(12), CK => n35, RESET => n8, Q => Q(12));
   D_I_13 : FD_1737 port map( D => d(13), CK => n35, RESET => n8, Q => Q(13));
   D_I_14 : FD_1736 port map( D => d(14), CK => n35, RESET => n8, Q => Q(14));
   D_I_15 : FD_1735 port map( D => d(15), CK => n35, RESET => n8, Q => Q(15));
   D_I_16 : FD_1734 port map( D => d(16), CK => n35, RESET => n8, Q => Q(16));
   D_I_17 : FD_1733 port map( D => d(17), CK => n35, RESET => n8, Q => Q(17));
   D_I_18 : FD_1732 port map( D => d(18), CK => n35, RESET => n8, Q => Q(18));
   D_I_19 : FD_1731 port map( D => d(19), CK => n35, RESET => n8, Q => Q(19));
   D_I_20 : FD_1730 port map( D => d(20), CK => n35, RESET => n8, Q => Q(20));
   D_I_21 : FD_1729 port map( D => d(21), CK => n35, RESET => n8, Q => Q(21));
   D_I_22 : FD_1728 port map( D => d(22), CK => n36, RESET => n8, Q => Q(22));
   D_I_23 : FD_1727 port map( D => d(23), CK => n36, RESET => n8, Q => Q(23));
   D_I_24 : FD_1726 port map( D => d(24), CK => n36, RESET => n9, Q => Q(24));
   D_I_25 : FD_1725 port map( D => d(25), CK => n36, RESET => n9, Q => Q(25));
   D_I_26 : FD_1724 port map( D => d(26), CK => n36, RESET => n9, Q => Q(26));
   D_I_27 : FD_1723 port map( D => d(27), CK => n36, RESET => n9, Q => Q(27));
   D_I_28 : FD_1722 port map( D => d(28), CK => n36, RESET => n9, Q => Q(28));
   D_I_29 : FD_1721 port map( D => d(29), CK => n36, RESET => n9, Q => Q(29));
   D_I_30 : FD_1720 port map( D => d(30), CK => n36, RESET => n9, Q => Q(30));
   D_I_31 : FD_1719 port map( D => d(31), CK => n36, RESET => n9, Q => Q(31));
   D_I_32 : FD_1718 port map( D => d(32), CK => n36, RESET => n9, Q => Q(32));
   D_I_33 : FD_1717 port map( D => d(33), CK => n37, RESET => n9, Q => Q(33));
   D_I_34 : FD_1716 port map( D => d(34), CK => n37, RESET => n9, Q => Q(34));
   D_I_35 : FD_1715 port map( D => d(35), CK => n37, RESET => n9, Q => Q(35));
   D_I_36 : FD_1714 port map( D => d(36), CK => n37, RESET => n10, Q => Q(36));
   D_I_37 : FD_1713 port map( D => d(37), CK => n37, RESET => n10, Q => Q(37));
   D_I_38 : FD_1712 port map( D => d(38), CK => n37, RESET => n10, Q => Q(38));
   D_I_39 : FD_1711 port map( D => d(39), CK => n37, RESET => n10, Q => Q(39));
   D_I_40 : FD_1710 port map( D => d(40), CK => n37, RESET => n10, Q => Q(40));
   D_I_41 : FD_1709 port map( D => d(41), CK => n37, RESET => n10, Q => Q(41));
   D_I_42 : FD_1708 port map( D => d(42), CK => n37, RESET => n10, Q => Q(42));
   D_I_43 : FD_1707 port map( D => d(43), CK => n37, RESET => n10, Q => Q(43));
   D_I_44 : FD_1706 port map( D => d(44), CK => n38, RESET => n10, Q => Q(44));
   D_I_45 : FD_1705 port map( D => d(45), CK => n38, RESET => n10, Q => Q(45));
   D_I_46 : FD_1704 port map( D => d(46), CK => n38, RESET => n10, Q => Q(46));
   D_I_47 : FD_1703 port map( D => d(47), CK => n38, RESET => n10, Q => Q(47));
   D_I_48 : FD_1702 port map( D => d(48), CK => n38, RESET => n11, Q => Q(48));
   D_I_49 : FD_1701 port map( D => d(49), CK => n38, RESET => n11, Q => Q(49));
   D_I_50 : FD_1700 port map( D => d(50), CK => n38, RESET => n11, Q => Q(50));
   D_I_51 : FD_1699 port map( D => d(51), CK => n38, RESET => n11, Q => Q(51));
   D_I_52 : FD_1698 port map( D => d(52), CK => n38, RESET => n11, Q => Q(52));
   D_I_53 : FD_1697 port map( D => d(53), CK => n38, RESET => n11, Q => Q(53));
   D_I_54 : FD_1696 port map( D => d(54), CK => n38, RESET => n11, Q => Q(54));
   D_I_55 : FD_1695 port map( D => d(55), CK => n39, RESET => n11, Q => Q(55));
   D_I_56 : FD_1694 port map( D => d(56), CK => n39, RESET => n11, Q => Q(56));
   D_I_57 : FD_1693 port map( D => d(57), CK => n39, RESET => n11, Q => Q(57));
   D_I_58 : FD_1692 port map( D => d(58), CK => n39, RESET => n11, Q => Q(58));
   D_I_59 : FD_1691 port map( D => d(59), CK => n39, RESET => n11, Q => Q(59));
   D_I_60 : FD_1690 port map( D => d(60), CK => n39, RESET => n12, Q => Q(60));
   D_I_61 : FD_1689 port map( D => d(61), CK => n39, RESET => n12, Q => Q(61));
   D_I_62 : FD_1688 port map( D => d(62), CK => n39, RESET => n12, Q => Q(62));
   D_I_63 : FD_1687 port map( D => d(63), CK => n39, RESET => n12, Q => Q(63));
   D_I_64 : FD_1686 port map( D => d(64), CK => n39, RESET => n12, Q => Q(64));
   D_I_65 : FD_1685 port map( D => d(65), CK => n39, RESET => n12, Q => Q(65));
   D_I_66 : FD_1684 port map( D => d(66), CK => n40, RESET => n12, Q => Q(66));
   D_I_67 : FD_1683 port map( D => d(67), CK => n40, RESET => n12, Q => Q(67));
   D_I_68 : FD_1682 port map( D => d(68), CK => n40, RESET => n12, Q => Q(68));
   D_I_69 : FD_1681 port map( D => d(69), CK => n40, RESET => n12, Q => Q(69));
   D_I_70 : FD_1680 port map( D => d(70), CK => n40, RESET => n12, Q => Q(70));
   D_I_71 : FD_1679 port map( D => d(71), CK => n40, RESET => n12, Q => Q(71));
   D_I_72 : FD_1678 port map( D => d(72), CK => n40, RESET => n13, Q => Q(72));
   D_I_73 : FD_1677 port map( D => d(73), CK => n40, RESET => n13, Q => Q(73));
   D_I_74 : FD_1676 port map( D => d(74), CK => n40, RESET => n13, Q => Q(74));
   D_I_75 : FD_1675 port map( D => d(75), CK => n40, RESET => n13, Q => Q(75));
   D_I_76 : FD_1674 port map( D => d(76), CK => n40, RESET => n13, Q => Q(76));
   D_I_77 : FD_1673 port map( D => d(77), CK => n41, RESET => n13, Q => Q(77));
   D_I_78 : FD_1672 port map( D => d(78), CK => n41, RESET => n13, Q => Q(78));
   D_I_79 : FD_1671 port map( D => d(79), CK => n41, RESET => n13, Q => Q(79));
   D_I_80 : FD_1670 port map( D => d(80), CK => n41, RESET => n13, Q => Q(80));
   D_I_81 : FD_1669 port map( D => d(81), CK => n41, RESET => n13, Q => Q(81));
   D_I_82 : FD_1668 port map( D => d(82), CK => n41, RESET => n13, Q => Q(82));
   D_I_83 : FD_1667 port map( D => d(83), CK => n41, RESET => n13, Q => Q(83));
   D_I_84 : FD_1666 port map( D => d(84), CK => n41, RESET => n14, Q => Q(84));
   D_I_85 : FD_1665 port map( D => d(85), CK => n41, RESET => n14, Q => Q(85));
   D_I_86 : FD_1664 port map( D => d(86), CK => n41, RESET => n14, Q => Q(86));
   D_I_87 : FD_1663 port map( D => d(87), CK => n41, RESET => n14, Q => Q(87));
   D_I_88 : FD_1662 port map( D => d(88), CK => n42, RESET => n14, Q => Q(88));
   D_I_89 : FD_1661 port map( D => d(89), CK => n42, RESET => n14, Q => Q(89));
   D_I_90 : FD_1660 port map( D => d(90), CK => n42, RESET => n14, Q => Q(90));
   D_I_91 : FD_1659 port map( D => d(91), CK => n42, RESET => n14, Q => Q(91));
   D_I_92 : FD_1658 port map( D => d(92), CK => n42, RESET => n14, Q => Q(92));
   D_I_93 : FD_1657 port map( D => d(93), CK => n42, RESET => n14, Q => Q(93));
   D_I_94 : FD_1656 port map( D => d(94), CK => n42, RESET => n14, Q => Q(94));
   D_I_95 : FD_1655 port map( D => d(95), CK => n42, RESET => n14, Q => Q(95));
   D_I_96 : FD_1654 port map( D => d(96), CK => n42, RESET => n15, Q => Q(96));
   D_I_97 : FD_1653 port map( D => d(97), CK => n42, RESET => n15, Q => Q(97));
   D_I_98 : FD_1652 port map( D => d(98), CK => n42, RESET => n15, Q => Q(98));
   D_I_99 : FD_1651 port map( D => d(99), CK => n43, RESET => n15, Q => Q(99));
   D_I_100 : FD_1650 port map( D => d(100), CK => n43, RESET => n15, Q => 
                           Q(100));
   D_I_101 : FD_1649 port map( D => d(101), CK => n43, RESET => n15, Q => 
                           Q(101));
   D_I_102 : FD_1648 port map( D => d(102), CK => n43, RESET => n15, Q => 
                           Q(102));
   D_I_103 : FD_1647 port map( D => d(103), CK => n43, RESET => n15, Q => 
                           Q(103));
   D_I_104 : FD_1646 port map( D => d(104), CK => n43, RESET => n15, Q => 
                           Q(104));
   D_I_105 : FD_1645 port map( D => d(105), CK => n43, RESET => n15, Q => 
                           Q(105));
   D_I_106 : FD_1644 port map( D => d(106), CK => n43, RESET => n15, Q => 
                           Q(106));
   D_I_107 : FD_1643 port map( D => d(107), CK => n43, RESET => n15, Q => 
                           Q(107));
   D_I_108 : FD_1642 port map( D => d(108), CK => n43, RESET => n16, Q => 
                           Q(108));
   D_I_109 : FD_1641 port map( D => d(109), CK => n43, RESET => n16, Q => 
                           Q(109));
   D_I_110 : FD_1640 port map( D => d(110), CK => n44, RESET => n16, Q => 
                           Q(110));
   D_I_111 : FD_1639 port map( D => d(111), CK => n44, RESET => n16, Q => 
                           Q(111));
   D_I_112 : FD_1638 port map( D => d(112), CK => n44, RESET => n16, Q => 
                           Q(112));
   D_I_113 : FD_1637 port map( D => d(113), CK => n44, RESET => n16, Q => 
                           Q(113));
   D_I_114 : FD_1636 port map( D => d(114), CK => n44, RESET => n16, Q => 
                           Q(114));
   D_I_115 : FD_1635 port map( D => d(115), CK => n44, RESET => n16, Q => 
                           Q(115));
   D_I_116 : FD_1634 port map( D => d(116), CK => n44, RESET => n16, Q => 
                           Q(116));
   D_I_117 : FD_1633 port map( D => d(117), CK => n44, RESET => n16, Q => 
                           Q(117));
   D_I_118 : FD_1632 port map( D => d(118), CK => n44, RESET => n16, Q => 
                           Q(118));
   D_I_119 : FD_1631 port map( D => d(119), CK => n44, RESET => n16, Q => 
                           Q(119));
   D_I_120 : FD_1630 port map( D => d(120), CK => n44, RESET => n17, Q => 
                           Q(120));
   D_I_121 : FD_1629 port map( D => d(121), CK => n45, RESET => n17, Q => 
                           Q(121));
   D_I_122 : FD_1628 port map( D => d(122), CK => n45, RESET => n17, Q => 
                           Q(122));
   D_I_123 : FD_1627 port map( D => d(123), CK => n45, RESET => n17, Q => 
                           Q(123));
   D_I_124 : FD_1626 port map( D => d(124), CK => n45, RESET => n17, Q => 
                           Q(124));
   D_I_125 : FD_1625 port map( D => d(125), CK => n45, RESET => n17, Q => 
                           Q(125));
   D_I_126 : FD_1624 port map( D => d(126), CK => n45, RESET => n17, Q => 
                           Q(126));
   D_I_127 : FD_1623 port map( D => d(127), CK => n45, RESET => n17, Q => 
                           Q(127));
   D_I_128 : FD_1622 port map( D => d(128), CK => n45, RESET => n17, Q => 
                           Q(128));
   D_I_129 : FD_1621 port map( D => d(129), CK => n45, RESET => n17, Q => 
                           Q(129));
   D_I_130 : FD_1620 port map( D => d(130), CK => n45, RESET => n17, Q => 
                           Q(130));
   D_I_131 : FD_1619 port map( D => d(131), CK => n45, RESET => n17, Q => 
                           Q(131));
   D_I_132 : FD_1618 port map( D => d(132), CK => n46, RESET => n18, Q => 
                           Q(132));
   D_I_133 : FD_1617 port map( D => d(133), CK => n46, RESET => n18, Q => 
                           Q(133));
   D_I_134 : FD_1616 port map( D => d(134), CK => n46, RESET => n18, Q => 
                           Q(134));
   D_I_135 : FD_1615 port map( D => d(135), CK => n46, RESET => n18, Q => 
                           Q(135));
   D_I_136 : FD_1614 port map( D => d(136), CK => n46, RESET => n18, Q => 
                           Q(136));
   D_I_137 : FD_1613 port map( D => d(137), CK => n46, RESET => n18, Q => 
                           Q(137));
   D_I_138 : FD_1612 port map( D => d(138), CK => n46, RESET => n18, Q => 
                           Q(138));
   D_I_139 : FD_1611 port map( D => d(139), CK => n46, RESET => n18, Q => 
                           Q(139));
   D_I_140 : FD_1610 port map( D => d(140), CK => n46, RESET => n18, Q => 
                           Q(140));
   D_I_141 : FD_1609 port map( D => d(141), CK => n46, RESET => n18, Q => 
                           Q(141));
   D_I_142 : FD_1608 port map( D => d(142), CK => n46, RESET => n18, Q => 
                           Q(142));
   D_I_143 : FD_1607 port map( D => d(143), CK => n47, RESET => n18, Q => 
                           Q(143));
   D_I_144 : FD_1606 port map( D => d(144), CK => n47, RESET => n19, Q => 
                           Q(144));
   D_I_145 : FD_1605 port map( D => d(145), CK => n47, RESET => n19, Q => 
                           Q(145));
   D_I_146 : FD_1604 port map( D => d(146), CK => n47, RESET => n19, Q => 
                           Q(146));
   D_I_147 : FD_1603 port map( D => d(147), CK => n47, RESET => n19, Q => 
                           Q(147));
   D_I_148 : FD_1602 port map( D => d(148), CK => n47, RESET => n19, Q => 
                           Q(148));
   D_I_149 : FD_1601 port map( D => d(149), CK => n47, RESET => n19, Q => 
                           Q(149));
   D_I_150 : FD_1600 port map( D => d(150), CK => n47, RESET => n19, Q => 
                           Q(150));
   D_I_151 : FD_1599 port map( D => d(151), CK => n47, RESET => n19, Q => 
                           Q(151));
   D_I_152 : FD_1598 port map( D => d(152), CK => n47, RESET => n19, Q => 
                           Q(152));
   D_I_153 : FD_1597 port map( D => d(153), CK => n47, RESET => n19, Q => 
                           Q(153));
   D_I_154 : FD_1596 port map( D => d(154), CK => n48, RESET => n19, Q => 
                           Q(154));
   D_I_155 : FD_1595 port map( D => d(155), CK => n48, RESET => n19, Q => 
                           Q(155));
   D_I_156 : FD_1594 port map( D => d(156), CK => n48, RESET => n20, Q => 
                           Q(156));
   D_I_157 : FD_1593 port map( D => d(157), CK => n48, RESET => n20, Q => 
                           Q(157));
   D_I_158 : FD_1592 port map( D => d(158), CK => n48, RESET => n20, Q => 
                           Q(158));
   D_I_159 : FD_1591 port map( D => d(159), CK => n48, RESET => n20, Q => 
                           Q(159));
   D_I_160 : FD_1590 port map( D => d(160), CK => n48, RESET => n20, Q => 
                           Q(160));
   D_I_161 : FD_1589 port map( D => d(161), CK => n48, RESET => n20, Q => 
                           Q(161));
   D_I_162 : FD_1588 port map( D => d(162), CK => n48, RESET => n20, Q => 
                           Q(162));
   D_I_163 : FD_1587 port map( D => d(163), CK => n48, RESET => n20, Q => 
                           Q(163));
   D_I_164 : FD_1586 port map( D => d(164), CK => n48, RESET => n20, Q => 
                           Q(164));
   D_I_165 : FD_1585 port map( D => d(165), CK => n49, RESET => n20, Q => 
                           Q(165));
   D_I_166 : FD_1584 port map( D => d(166), CK => n49, RESET => n20, Q => 
                           Q(166));
   D_I_167 : FD_1583 port map( D => d(167), CK => n49, RESET => n20, Q => 
                           Q(167));
   D_I_168 : FD_1582 port map( D => d(168), CK => n49, RESET => n21, Q => 
                           Q(168));
   D_I_169 : FD_1581 port map( D => d(169), CK => n49, RESET => n21, Q => 
                           Q(169));
   D_I_170 : FD_1580 port map( D => d(170), CK => n49, RESET => n21, Q => 
                           Q(170));
   D_I_171 : FD_1579 port map( D => d(171), CK => n49, RESET => n21, Q => 
                           Q(171));
   D_I_172 : FD_1578 port map( D => d(172), CK => n49, RESET => n21, Q => 
                           Q(172));
   D_I_173 : FD_1577 port map( D => d(173), CK => n49, RESET => n21, Q => 
                           Q(173));
   D_I_174 : FD_1576 port map( D => d(174), CK => n49, RESET => n21, Q => 
                           Q(174));
   D_I_175 : FD_1575 port map( D => d(175), CK => n49, RESET => n21, Q => 
                           Q(175));
   D_I_176 : FD_1574 port map( D => d(176), CK => n50, RESET => n21, Q => 
                           Q(176));
   D_I_177 : FD_1573 port map( D => d(177), CK => n50, RESET => n21, Q => 
                           Q(177));
   D_I_178 : FD_1572 port map( D => d(178), CK => n50, RESET => n21, Q => 
                           Q(178));
   D_I_179 : FD_1571 port map( D => d(179), CK => n50, RESET => n21, Q => 
                           Q(179));
   D_I_180 : FD_1570 port map( D => d(180), CK => n50, RESET => n22, Q => 
                           Q(180));
   D_I_181 : FD_1569 port map( D => d(181), CK => n50, RESET => n22, Q => 
                           Q(181));
   D_I_182 : FD_1568 port map( D => d(182), CK => n50, RESET => n22, Q => 
                           Q(182));
   D_I_183 : FD_1567 port map( D => d(183), CK => n50, RESET => n22, Q => 
                           Q(183));
   D_I_184 : FD_1566 port map( D => d(184), CK => n50, RESET => n22, Q => 
                           Q(184));
   D_I_185 : FD_1565 port map( D => d(185), CK => n50, RESET => n22, Q => 
                           Q(185));
   D_I_186 : FD_1564 port map( D => d(186), CK => n50, RESET => n22, Q => 
                           Q(186));
   D_I_187 : FD_1563 port map( D => d(187), CK => n51, RESET => n22, Q => 
                           Q(187));
   D_I_188 : FD_1562 port map( D => d(188), CK => n51, RESET => n22, Q => 
                           Q(188));
   D_I_189 : FD_1561 port map( D => d(189), CK => n51, RESET => n22, Q => 
                           Q(189));
   D_I_190 : FD_1560 port map( D => d(190), CK => n51, RESET => n22, Q => 
                           Q(190));
   D_I_191 : FD_1559 port map( D => d(191), CK => n51, RESET => n22, Q => 
                           Q(191));
   D_I_192 : FD_1558 port map( D => d(192), CK => n51, RESET => n23, Q => 
                           Q(192));
   D_I_193 : FD_1557 port map( D => d(193), CK => n51, RESET => n23, Q => 
                           Q(193));
   D_I_194 : FD_1556 port map( D => d(194), CK => n51, RESET => n23, Q => 
                           Q(194));
   D_I_195 : FD_1555 port map( D => d(195), CK => n51, RESET => n23, Q => 
                           Q(195));
   D_I_196 : FD_1554 port map( D => d(196), CK => n51, RESET => n23, Q => 
                           Q(196));
   D_I_197 : FD_1553 port map( D => d(197), CK => n51, RESET => n23, Q => 
                           Q(197));
   D_I_198 : FD_1552 port map( D => d(198), CK => n52, RESET => n23, Q => 
                           Q(198));
   D_I_199 : FD_1551 port map( D => d(199), CK => n52, RESET => n23, Q => 
                           Q(199));
   D_I_200 : FD_1550 port map( D => d(200), CK => n52, RESET => n23, Q => 
                           Q(200));
   D_I_201 : FD_1549 port map( D => d(201), CK => n52, RESET => n23, Q => 
                           Q(201));
   D_I_202 : FD_1548 port map( D => d(202), CK => n52, RESET => n23, Q => 
                           Q(202));
   D_I_203 : FD_1547 port map( D => d(203), CK => n52, RESET => n23, Q => 
                           Q(203));
   D_I_204 : FD_1546 port map( D => d(204), CK => n52, RESET => n24, Q => 
                           Q(204));
   D_I_205 : FD_1545 port map( D => d(205), CK => n52, RESET => n24, Q => 
                           Q(205));
   D_I_206 : FD_1544 port map( D => d(206), CK => n52, RESET => n24, Q => 
                           Q(206));
   D_I_207 : FD_1543 port map( D => d(207), CK => n52, RESET => n24, Q => 
                           Q(207));
   D_I_208 : FD_1542 port map( D => d(208), CK => n52, RESET => n24, Q => 
                           Q(208));
   D_I_209 : FD_1541 port map( D => d(209), CK => n53, RESET => n24, Q => 
                           Q(209));
   D_I_210 : FD_1540 port map( D => d(210), CK => n53, RESET => n24, Q => 
                           Q(210));
   D_I_211 : FD_1539 port map( D => d(211), CK => n53, RESET => n24, Q => 
                           Q(211));
   D_I_212 : FD_1538 port map( D => d(212), CK => n53, RESET => n24, Q => 
                           Q(212));
   D_I_213 : FD_1537 port map( D => d(213), CK => n53, RESET => n24, Q => 
                           Q(213));
   D_I_214 : FD_1536 port map( D => d(214), CK => n53, RESET => n24, Q => 
                           Q(214));
   D_I_215 : FD_1535 port map( D => d(215), CK => n53, RESET => n24, Q => 
                           Q(215));
   D_I_216 : FD_1534 port map( D => d(216), CK => n53, RESET => n25, Q => 
                           Q(216));
   D_I_217 : FD_1533 port map( D => d(217), CK => n53, RESET => n25, Q => 
                           Q(217));
   D_I_218 : FD_1532 port map( D => d(218), CK => n53, RESET => n25, Q => 
                           Q(218));
   D_I_219 : FD_1531 port map( D => d(219), CK => n53, RESET => n25, Q => 
                           Q(219));
   D_I_220 : FD_1530 port map( D => d(220), CK => n54, RESET => n25, Q => 
                           Q(220));
   D_I_221 : FD_1529 port map( D => d(221), CK => n54, RESET => n25, Q => 
                           Q(221));
   D_I_222 : FD_1528 port map( D => d(222), CK => n54, RESET => n25, Q => 
                           Q(222));
   D_I_223 : FD_1527 port map( D => d(223), CK => n54, RESET => n25, Q => 
                           Q(223));
   D_I_224 : FD_1526 port map( D => d(224), CK => n54, RESET => n25, Q => 
                           Q(224));
   D_I_225 : FD_1525 port map( D => d(225), CK => n54, RESET => n25, Q => 
                           Q(225));
   D_I_226 : FD_1524 port map( D => d(226), CK => n54, RESET => n25, Q => 
                           Q(226));
   D_I_227 : FD_1523 port map( D => d(227), CK => n54, RESET => n25, Q => 
                           Q(227));
   D_I_228 : FD_1522 port map( D => d(228), CK => n54, RESET => n26, Q => 
                           Q(228));
   D_I_229 : FD_1521 port map( D => d(229), CK => n54, RESET => n26, Q => 
                           Q(229));
   D_I_230 : FD_1520 port map( D => d(230), CK => n54, RESET => n26, Q => 
                           Q(230));
   D_I_231 : FD_1519 port map( D => d(231), CK => n55, RESET => n26, Q => 
                           Q(231));
   D_I_232 : FD_1518 port map( D => d(232), CK => n55, RESET => n26, Q => 
                           Q(232));
   D_I_233 : FD_1517 port map( D => d(233), CK => n55, RESET => n26, Q => 
                           Q(233));
   D_I_234 : FD_1516 port map( D => d(234), CK => n55, RESET => n26, Q => 
                           Q(234));
   D_I_235 : FD_1515 port map( D => d(235), CK => n55, RESET => n26, Q => 
                           Q(235));
   D_I_236 : FD_1514 port map( D => d(236), CK => n55, RESET => n26, Q => 
                           Q(236));
   D_I_237 : FD_1513 port map( D => d(237), CK => n55, RESET => n26, Q => 
                           Q(237));
   D_I_238 : FD_1512 port map( D => d(238), CK => n55, RESET => n26, Q => 
                           Q(238));
   D_I_239 : FD_1511 port map( D => d(239), CK => n55, RESET => n26, Q => 
                           Q(239));
   D_I_240 : FD_1510 port map( D => d(240), CK => n55, RESET => n27, Q => 
                           Q(240));
   D_I_241 : FD_1509 port map( D => d(241), CK => n55, RESET => n27, Q => 
                           Q(241));
   D_I_242 : FD_1508 port map( D => d(242), CK => n56, RESET => n27, Q => 
                           Q(242));
   D_I_243 : FD_1507 port map( D => d(243), CK => n56, RESET => n27, Q => 
                           Q(243));
   D_I_244 : FD_1506 port map( D => d(244), CK => n56, RESET => n27, Q => 
                           Q(244));
   D_I_245 : FD_1505 port map( D => d(245), CK => n56, RESET => n27, Q => 
                           Q(245));
   D_I_246 : FD_1504 port map( D => d(246), CK => n56, RESET => n27, Q => 
                           Q(246));
   D_I_247 : FD_1503 port map( D => d(247), CK => n56, RESET => n27, Q => 
                           Q(247));
   D_I_248 : FD_1502 port map( D => d(248), CK => n56, RESET => n27, Q => 
                           Q(248));
   U1 : BUF_X1 port map( A => n6, Z => n1);
   U2 : BUF_X1 port map( A => n6, Z => n2);
   U3 : BUF_X1 port map( A => n5, Z => n3);
   U4 : BUF_X1 port map( A => n5, Z => n4);
   U5 : BUF_X1 port map( A => n33, Z => n28);
   U6 : BUF_X1 port map( A => n33, Z => n29);
   U7 : BUF_X1 port map( A => n32, Z => n30);
   U8 : BUF_X1 port map( A => n32, Z => n31);
   U9 : BUF_X1 port map( A => reset, Z => n6);
   U10 : BUF_X1 port map( A => reset, Z => n5);
   U11 : BUF_X1 port map( A => clk, Z => n33);
   U12 : BUF_X1 port map( A => clk, Z => n32);
   U13 : CLKBUF_X1 port map( A => n1, Z => n7);
   U14 : CLKBUF_X1 port map( A => n1, Z => n8);
   U15 : CLKBUF_X1 port map( A => n1, Z => n9);
   U16 : CLKBUF_X1 port map( A => n1, Z => n10);
   U17 : CLKBUF_X1 port map( A => n1, Z => n11);
   U18 : CLKBUF_X1 port map( A => n1, Z => n12);
   U19 : CLKBUF_X1 port map( A => n2, Z => n13);
   U20 : CLKBUF_X1 port map( A => n2, Z => n14);
   U21 : CLKBUF_X1 port map( A => n2, Z => n15);
   U22 : CLKBUF_X1 port map( A => n2, Z => n16);
   U23 : CLKBUF_X1 port map( A => n2, Z => n17);
   U24 : CLKBUF_X1 port map( A => n2, Z => n18);
   U25 : CLKBUF_X1 port map( A => n3, Z => n19);
   U26 : CLKBUF_X1 port map( A => n3, Z => n20);
   U27 : CLKBUF_X1 port map( A => n3, Z => n21);
   U28 : CLKBUF_X1 port map( A => n3, Z => n22);
   U29 : CLKBUF_X1 port map( A => n3, Z => n23);
   U30 : CLKBUF_X1 port map( A => n3, Z => n24);
   U31 : CLKBUF_X1 port map( A => n4, Z => n25);
   U32 : CLKBUF_X1 port map( A => n4, Z => n26);
   U33 : CLKBUF_X1 port map( A => n4, Z => n27);
   U34 : CLKBUF_X1 port map( A => n28, Z => n34);
   U35 : CLKBUF_X1 port map( A => n28, Z => n35);
   U36 : CLKBUF_X1 port map( A => n28, Z => n36);
   U37 : CLKBUF_X1 port map( A => n28, Z => n37);
   U38 : CLKBUF_X1 port map( A => n28, Z => n38);
   U39 : CLKBUF_X1 port map( A => n28, Z => n39);
   U40 : CLKBUF_X1 port map( A => n29, Z => n40);
   U41 : CLKBUF_X1 port map( A => n29, Z => n41);
   U42 : CLKBUF_X1 port map( A => n29, Z => n42);
   U43 : CLKBUF_X1 port map( A => n29, Z => n43);
   U44 : CLKBUF_X1 port map( A => n29, Z => n44);
   U45 : CLKBUF_X1 port map( A => n29, Z => n45);
   U46 : CLKBUF_X1 port map( A => n30, Z => n46);
   U47 : CLKBUF_X1 port map( A => n30, Z => n47);
   U48 : CLKBUF_X1 port map( A => n30, Z => n48);
   U49 : CLKBUF_X1 port map( A => n30, Z => n49);
   U50 : CLKBUF_X1 port map( A => n30, Z => n50);
   U51 : CLKBUF_X1 port map( A => n30, Z => n51);
   U52 : CLKBUF_X1 port map( A => n31, Z => n52);
   U53 : CLKBUF_X1 port map( A => n31, Z => n53);
   U54 : CLKBUF_X1 port map( A => n31, Z => n54);
   U55 : CLKBUF_X1 port map( A => n31, Z => n55);
   U56 : CLKBUF_X1 port map( A => n31, Z => n56);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity adder_NBIT19 is

   port( a, b : in std_logic_vector (18 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (19 downto 0));

end adder_NBIT19;

architecture SYN_beh of adder_NBIT19 is

   component adder_NBIT19_DW01_add_0
      port( A, B : in std_logic_vector (19 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (19 downto 0);  CO : out std_logic);
   end component;
   
   signal n_3355 : std_logic;

begin
   
   add_1_root_add_21_2 : adder_NBIT19_DW01_add_0 port map( A(19) => a(18), 
                           A(18) => a(18), A(17) => a(17), A(16) => a(16), 
                           A(15) => a(15), A(14) => a(14), A(13) => a(13), 
                           A(12) => a(12), A(11) => a(11), A(10) => a(10), A(9)
                           => a(9), A(8) => a(8), A(7) => a(7), A(6) => a(6), 
                           A(5) => a(5), A(4) => a(4), A(3) => a(3), A(2) => 
                           a(2), A(1) => a(1), A(0) => a(0), B(19) => b(18), 
                           B(18) => b(18), B(17) => b(17), B(16) => b(16), 
                           B(15) => b(15), B(14) => b(14), B(13) => b(13), 
                           B(12) => b(12), B(11) => b(11), B(10) => b(10), B(9)
                           => b(9), B(8) => b(8), B(7) => b(7), B(6) => b(6), 
                           B(5) => b(5), B(4) => b(4), B(3) => b(3), B(2) => 
                           b(2), B(1) => b(1), B(0) => b(0), CI => cin, SUM(19)
                           => s(19), SUM(18) => s(18), SUM(17) => s(17), 
                           SUM(16) => s(16), SUM(15) => s(15), SUM(14) => s(14)
                           , SUM(13) => s(13), SUM(12) => s(12), SUM(11) => 
                           s(11), SUM(10) => s(10), SUM(9) => s(9), SUM(8) => 
                           s(8), SUM(7) => s(7), SUM(6) => s(6), SUM(5) => s(5)
                           , SUM(4) => s(4), SUM(3) => s(3), SUM(2) => s(2), 
                           SUM(1) => s(1), SUM(0) => s(0), CO => n_3355);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N19_Z3 is

   port( inputs : in std_logic_vector (0 to 151);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (18 downto 0));

end MUX_zbit_nbit_N19_Z3;

architecture SYN_beh of MUX_zbit_nbit_N19_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, 
      N146, N147, N148, N149, N150, N151, N152, N153, n4, n1, n2, n3, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90 : std_logic;

begin
   
   Y_reg_18_inst : DLH_X1 port map( G => n4, D => N153, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n4, D => N152, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N151, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N150, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N149, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N148, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N147, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N146, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N145, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N144, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N143, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N142, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N141, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N140, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N139, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N138, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N137, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N136, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N135, Q => Y(0));
   n4 <= '1';
   U3 : OR4_X1 port map( A1 => n9, A2 => n10, A3 => n8, A4 => n87, ZN => n7);
   U4 : INV_X1 port map( A => n7, ZN => n1);
   U5 : NOR3_X4 port map( A1 => n88, A2 => SEL(1), A3 => n90, ZN => n12);
   U6 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(1), A3 => n88, ZN => n14);
   U7 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(2), A3 => n89, ZN => n11);
   U8 : NOR3_X4 port map( A1 => n90, A2 => n88, A3 => n89, ZN => n13);
   U9 : NOR3_X4 port map( A1 => n90, A2 => SEL(2), A3 => n89, ZN => n10);
   U10 : NOR3_X4 port map( A1 => n88, A2 => SEL(0), A3 => n89, ZN => n8);
   U11 : NOR3_X4 port map( A1 => SEL(1), A2 => SEL(2), A3 => n90, ZN => n9);
   U12 : NAND4_X1 port map( A1 => n2, A2 => n3, A3 => n5, A4 => n6, ZN => N153)
                           ;
   U13 : AOI22_X1 port map( A1 => inputs(0), A2 => n1, B1 => inputs(114), B2 =>
                           n8, ZN => n6);
   U14 : AOI22_X1 port map( A1 => inputs(19), A2 => n9, B1 => inputs(57), B2 =>
                           n10, ZN => n5);
   U15 : AOI22_X1 port map( A1 => inputs(38), A2 => n11, B1 => inputs(95), B2 
                           => n12, ZN => n3);
   U16 : AOI22_X1 port map( A1 => inputs(133), A2 => n13, B1 => inputs(76), B2 
                           => n14, ZN => n2);
   U17 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           N152);
   U18 : AOI22_X1 port map( A1 => inputs(1), A2 => n1, B1 => inputs(115), B2 =>
                           n8, ZN => n18);
   U19 : AOI22_X1 port map( A1 => inputs(20), A2 => n9, B1 => inputs(58), B2 =>
                           n10, ZN => n17);
   U20 : AOI22_X1 port map( A1 => inputs(39), A2 => n11, B1 => inputs(96), B2 
                           => n12, ZN => n16);
   U21 : AOI22_X1 port map( A1 => inputs(134), A2 => n13, B1 => inputs(77), B2 
                           => n14, ZN => n15);
   U22 : NAND4_X1 port map( A1 => n19, A2 => n20, A3 => n21, A4 => n22, ZN => 
                           N151);
   U23 : AOI22_X1 port map( A1 => inputs(2), A2 => n1, B1 => inputs(116), B2 =>
                           n8, ZN => n22);
   U24 : AOI22_X1 port map( A1 => inputs(21), A2 => n9, B1 => inputs(59), B2 =>
                           n10, ZN => n21);
   U25 : AOI22_X1 port map( A1 => inputs(40), A2 => n11, B1 => inputs(97), B2 
                           => n12, ZN => n20);
   U26 : AOI22_X1 port map( A1 => inputs(135), A2 => n13, B1 => inputs(78), B2 
                           => n14, ZN => n19);
   U27 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           N150);
   U28 : AOI22_X1 port map( A1 => inputs(3), A2 => n1, B1 => inputs(117), B2 =>
                           n8, ZN => n26);
   U29 : AOI22_X1 port map( A1 => inputs(22), A2 => n9, B1 => inputs(60), B2 =>
                           n10, ZN => n25);
   U30 : AOI22_X1 port map( A1 => inputs(41), A2 => n11, B1 => inputs(98), B2 
                           => n12, ZN => n24);
   U31 : AOI22_X1 port map( A1 => inputs(136), A2 => n13, B1 => inputs(79), B2 
                           => n14, ZN => n23);
   U32 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n30, ZN => 
                           N149);
   U33 : AOI22_X1 port map( A1 => inputs(4), A2 => n1, B1 => inputs(118), B2 =>
                           n8, ZN => n30);
   U34 : AOI22_X1 port map( A1 => inputs(23), A2 => n9, B1 => inputs(61), B2 =>
                           n10, ZN => n29);
   U35 : AOI22_X1 port map( A1 => inputs(42), A2 => n11, B1 => inputs(99), B2 
                           => n12, ZN => n28);
   U36 : AOI22_X1 port map( A1 => inputs(137), A2 => n13, B1 => inputs(80), B2 
                           => n14, ZN => n27);
   U37 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           N148);
   U38 : AOI22_X1 port map( A1 => inputs(5), A2 => n1, B1 => inputs(119), B2 =>
                           n8, ZN => n34);
   U39 : AOI22_X1 port map( A1 => inputs(24), A2 => n9, B1 => inputs(62), B2 =>
                           n10, ZN => n33);
   U40 : AOI22_X1 port map( A1 => inputs(43), A2 => n11, B1 => inputs(100), B2 
                           => n12, ZN => n32);
   U41 : AOI22_X1 port map( A1 => inputs(138), A2 => n13, B1 => inputs(81), B2 
                           => n14, ZN => n31);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           N147);
   U43 : AOI22_X1 port map( A1 => inputs(6), A2 => n1, B1 => inputs(120), B2 =>
                           n8, ZN => n38);
   U44 : AOI22_X1 port map( A1 => inputs(25), A2 => n9, B1 => inputs(63), B2 =>
                           n10, ZN => n37);
   U45 : AOI22_X1 port map( A1 => inputs(44), A2 => n11, B1 => inputs(101), B2 
                           => n12, ZN => n36);
   U46 : AOI22_X1 port map( A1 => inputs(139), A2 => n13, B1 => inputs(82), B2 
                           => n14, ZN => n35);
   U47 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           N146);
   U48 : AOI22_X1 port map( A1 => inputs(7), A2 => n1, B1 => inputs(121), B2 =>
                           n8, ZN => n42);
   U49 : AOI22_X1 port map( A1 => inputs(26), A2 => n9, B1 => inputs(64), B2 =>
                           n10, ZN => n41);
   U50 : AOI22_X1 port map( A1 => inputs(45), A2 => n11, B1 => inputs(102), B2 
                           => n12, ZN => n40);
   U51 : AOI22_X1 port map( A1 => inputs(140), A2 => n13, B1 => inputs(83), B2 
                           => n14, ZN => n39);
   U52 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           N145);
   U53 : AOI22_X1 port map( A1 => inputs(8), A2 => n1, B1 => inputs(122), B2 =>
                           n8, ZN => n46);
   U54 : AOI22_X1 port map( A1 => inputs(27), A2 => n9, B1 => inputs(65), B2 =>
                           n10, ZN => n45);
   U55 : AOI22_X1 port map( A1 => inputs(46), A2 => n11, B1 => inputs(103), B2 
                           => n12, ZN => n44);
   U56 : AOI22_X1 port map( A1 => inputs(141), A2 => n13, B1 => inputs(84), B2 
                           => n14, ZN => n43);
   U57 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           N144);
   U58 : AOI22_X1 port map( A1 => inputs(9), A2 => n1, B1 => inputs(123), B2 =>
                           n8, ZN => n50);
   U59 : AOI22_X1 port map( A1 => inputs(28), A2 => n9, B1 => inputs(66), B2 =>
                           n10, ZN => n49);
   U60 : AOI22_X1 port map( A1 => inputs(47), A2 => n11, B1 => inputs(104), B2 
                           => n12, ZN => n48);
   U61 : AOI22_X1 port map( A1 => inputs(142), A2 => n13, B1 => inputs(85), B2 
                           => n14, ZN => n47);
   U62 : NAND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           N143);
   U63 : AOI22_X1 port map( A1 => inputs(10), A2 => n1, B1 => inputs(124), B2 
                           => n8, ZN => n54);
   U64 : AOI22_X1 port map( A1 => inputs(29), A2 => n9, B1 => inputs(67), B2 =>
                           n10, ZN => n53);
   U65 : AOI22_X1 port map( A1 => inputs(48), A2 => n11, B1 => inputs(105), B2 
                           => n12, ZN => n52);
   U66 : AOI22_X1 port map( A1 => inputs(143), A2 => n13, B1 => inputs(86), B2 
                           => n14, ZN => n51);
   U67 : NAND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           N142);
   U68 : AOI22_X1 port map( A1 => inputs(11), A2 => n1, B1 => inputs(125), B2 
                           => n8, ZN => n58);
   U69 : AOI22_X1 port map( A1 => inputs(30), A2 => n9, B1 => inputs(68), B2 =>
                           n10, ZN => n57);
   U70 : AOI22_X1 port map( A1 => inputs(49), A2 => n11, B1 => inputs(106), B2 
                           => n12, ZN => n56);
   U71 : AOI22_X1 port map( A1 => inputs(144), A2 => n13, B1 => inputs(87), B2 
                           => n14, ZN => n55);
   U72 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           N141);
   U73 : AOI22_X1 port map( A1 => inputs(12), A2 => n1, B1 => inputs(126), B2 
                           => n8, ZN => n62);
   U74 : AOI22_X1 port map( A1 => inputs(31), A2 => n9, B1 => inputs(69), B2 =>
                           n10, ZN => n61);
   U75 : AOI22_X1 port map( A1 => inputs(50), A2 => n11, B1 => inputs(107), B2 
                           => n12, ZN => n60);
   U76 : AOI22_X1 port map( A1 => inputs(145), A2 => n13, B1 => inputs(88), B2 
                           => n14, ZN => n59);
   U77 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           N140);
   U78 : AOI22_X1 port map( A1 => inputs(13), A2 => n1, B1 => inputs(127), B2 
                           => n8, ZN => n66);
   U79 : AOI22_X1 port map( A1 => inputs(32), A2 => n9, B1 => inputs(70), B2 =>
                           n10, ZN => n65);
   U80 : AOI22_X1 port map( A1 => inputs(51), A2 => n11, B1 => inputs(108), B2 
                           => n12, ZN => n64);
   U81 : AOI22_X1 port map( A1 => inputs(146), A2 => n13, B1 => inputs(89), B2 
                           => n14, ZN => n63);
   U82 : NAND4_X1 port map( A1 => n67, A2 => n68, A3 => n69, A4 => n70, ZN => 
                           N139);
   U83 : AOI22_X1 port map( A1 => inputs(14), A2 => n1, B1 => inputs(128), B2 
                           => n8, ZN => n70);
   U84 : AOI22_X1 port map( A1 => inputs(33), A2 => n9, B1 => inputs(71), B2 =>
                           n10, ZN => n69);
   U85 : AOI22_X1 port map( A1 => inputs(52), A2 => n11, B1 => inputs(109), B2 
                           => n12, ZN => n68);
   U86 : AOI22_X1 port map( A1 => inputs(147), A2 => n13, B1 => inputs(90), B2 
                           => n14, ZN => n67);
   U87 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           N138);
   U88 : AOI22_X1 port map( A1 => inputs(15), A2 => n1, B1 => inputs(129), B2 
                           => n8, ZN => n74);
   U89 : AOI22_X1 port map( A1 => inputs(34), A2 => n9, B1 => inputs(72), B2 =>
                           n10, ZN => n73);
   U90 : AOI22_X1 port map( A1 => inputs(53), A2 => n11, B1 => inputs(110), B2 
                           => n12, ZN => n72);
   U91 : AOI22_X1 port map( A1 => inputs(148), A2 => n13, B1 => inputs(91), B2 
                           => n14, ZN => n71);
   U92 : NAND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           N137);
   U93 : AOI22_X1 port map( A1 => inputs(16), A2 => n1, B1 => inputs(130), B2 
                           => n8, ZN => n78);
   U94 : AOI22_X1 port map( A1 => inputs(35), A2 => n9, B1 => inputs(73), B2 =>
                           n10, ZN => n77);
   U95 : AOI22_X1 port map( A1 => inputs(54), A2 => n11, B1 => inputs(111), B2 
                           => n12, ZN => n76);
   U96 : AOI22_X1 port map( A1 => inputs(149), A2 => n13, B1 => inputs(92), B2 
                           => n14, ZN => n75);
   U97 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           N136);
   U98 : AOI22_X1 port map( A1 => inputs(17), A2 => n1, B1 => inputs(131), B2 
                           => n8, ZN => n82);
   U99 : AOI22_X1 port map( A1 => inputs(36), A2 => n9, B1 => inputs(74), B2 =>
                           n10, ZN => n81);
   U100 : AOI22_X1 port map( A1 => inputs(55), A2 => n11, B1 => inputs(112), B2
                           => n12, ZN => n80);
   U101 : AOI22_X1 port map( A1 => inputs(150), A2 => n13, B1 => inputs(93), B2
                           => n14, ZN => n79);
   U102 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           N135);
   U103 : AOI22_X1 port map( A1 => inputs(18), A2 => n1, B1 => inputs(132), B2 
                           => n8, ZN => n86);
   U104 : OR4_X1 port map( A1 => n14, A2 => n13, A3 => n12, A4 => n11, ZN => 
                           n87);
   U105 : AOI22_X1 port map( A1 => inputs(37), A2 => n9, B1 => inputs(75), B2 
                           => n10, ZN => n85);
   U106 : AOI22_X1 port map( A1 => inputs(56), A2 => n11, B1 => inputs(113), B2
                           => n12, ZN => n84);
   U107 : AOI22_X1 port map( A1 => inputs(151), A2 => n13, B1 => inputs(94), B2
                           => n14, ZN => n83);
   U108 : INV_X1 port map( A => SEL(1), ZN => n89);
   U109 : INV_X1 port map( A => SEL(2), ZN => n88);
   U111 : INV_X1 port map( A => SEL(0), ZN => n90);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N17_Z3 is

   port( inputs : in std_logic_vector (0 to 135);  SEL : in std_logic_vector (2
         downto 0);  Y : out std_logic_vector (16 downto 0));

end MUX_zbit_nbit_N17_Z3;

architecture SYN_beh of MUX_zbit_nbit_N17_Z3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, 
      N134, N135, N136, N137, N138, N139, n4, n1, n2, n3, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83 : std_logic;

begin
   
   Y_reg_16_inst : DLH_X1 port map( G => n4, D => N139, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n4, D => N138, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n4, D => N137, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n4, D => N136, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n4, D => N135, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n4, D => N134, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n4, D => N133, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n4, D => N132, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n4, D => N131, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n4, D => N130, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n4, D => N129, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n4, D => N128, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n4, D => N127, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n4, D => N126, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n4, D => N125, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n4, D => N124, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n4, D => N123, Q => Y(0));
   n4 <= '1';
   U3 : OR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n83, ZN => n1);
   U4 : OR3_X1 port map( A1 => n81, A2 => SEL(0), A3 => n82, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => n3);
   U6 : INV_X1 port map( A => n1, ZN => n5);
   U7 : NOR4_X4 port map( A1 => n5, A2 => n11, A3 => n3, A4 => n80, ZN => n10);
   U8 : NOR3_X4 port map( A1 => n83, A2 => SEL(2), A3 => n82, ZN => n11);
   U9 : NOR3_X4 port map( A1 => n81, A2 => SEL(1), A3 => n83, ZN => n13);
   U10 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(1), A3 => n81, ZN => n15);
   U11 : NOR3_X4 port map( A1 => SEL(0), A2 => SEL(2), A3 => n82, ZN => n12);
   U12 : NOR3_X4 port map( A1 => n83, A2 => n81, A3 => n82, ZN => n14);
   U13 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => N139)
                           ;
   U14 : AOI22_X1 port map( A1 => inputs(0), A2 => n10, B1 => inputs(102), B2 
                           => n3, ZN => n9);
   U15 : AOI22_X1 port map( A1 => inputs(17), A2 => n5, B1 => inputs(51), B2 =>
                           n11, ZN => n8);
   U16 : AOI22_X1 port map( A1 => inputs(34), A2 => n12, B1 => inputs(85), B2 
                           => n13, ZN => n7);
   U17 : AOI22_X1 port map( A1 => inputs(119), A2 => n14, B1 => inputs(68), B2 
                           => n15, ZN => n6);
   U18 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           N138);
   U19 : AOI22_X1 port map( A1 => inputs(1), A2 => n10, B1 => inputs(103), B2 
                           => n3, ZN => n19);
   U20 : AOI22_X1 port map( A1 => inputs(18), A2 => n5, B1 => inputs(52), B2 =>
                           n11, ZN => n18);
   U21 : AOI22_X1 port map( A1 => inputs(35), A2 => n12, B1 => inputs(86), B2 
                           => n13, ZN => n17);
   U22 : AOI22_X1 port map( A1 => inputs(120), A2 => n14, B1 => inputs(69), B2 
                           => n15, ZN => n16);
   U23 : NAND4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           N137);
   U24 : AOI22_X1 port map( A1 => inputs(2), A2 => n10, B1 => inputs(104), B2 
                           => n3, ZN => n23);
   U25 : AOI22_X1 port map( A1 => inputs(19), A2 => n5, B1 => inputs(53), B2 =>
                           n11, ZN => n22);
   U26 : AOI22_X1 port map( A1 => inputs(36), A2 => n12, B1 => inputs(87), B2 
                           => n13, ZN => n21);
   U27 : AOI22_X1 port map( A1 => inputs(121), A2 => n14, B1 => inputs(70), B2 
                           => n15, ZN => n20);
   U28 : NAND4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           N136);
   U29 : AOI22_X1 port map( A1 => inputs(3), A2 => n10, B1 => inputs(105), B2 
                           => n3, ZN => n27);
   U30 : AOI22_X1 port map( A1 => inputs(20), A2 => n5, B1 => inputs(54), B2 =>
                           n11, ZN => n26);
   U31 : AOI22_X1 port map( A1 => inputs(37), A2 => n12, B1 => inputs(88), B2 
                           => n13, ZN => n25);
   U32 : AOI22_X1 port map( A1 => inputs(122), A2 => n14, B1 => inputs(71), B2 
                           => n15, ZN => n24);
   U33 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           N135);
   U34 : AOI22_X1 port map( A1 => inputs(4), A2 => n10, B1 => inputs(106), B2 
                           => n3, ZN => n31);
   U35 : AOI22_X1 port map( A1 => inputs(21), A2 => n5, B1 => inputs(55), B2 =>
                           n11, ZN => n30);
   U36 : AOI22_X1 port map( A1 => inputs(38), A2 => n12, B1 => inputs(89), B2 
                           => n13, ZN => n29);
   U37 : AOI22_X1 port map( A1 => inputs(123), A2 => n14, B1 => inputs(72), B2 
                           => n15, ZN => n28);
   U38 : NAND4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => 
                           N134);
   U39 : AOI22_X1 port map( A1 => inputs(5), A2 => n10, B1 => inputs(107), B2 
                           => n3, ZN => n35);
   U40 : AOI22_X1 port map( A1 => inputs(22), A2 => n5, B1 => inputs(56), B2 =>
                           n11, ZN => n34);
   U41 : AOI22_X1 port map( A1 => inputs(39), A2 => n12, B1 => inputs(90), B2 
                           => n13, ZN => n33);
   U42 : AOI22_X1 port map( A1 => inputs(124), A2 => n14, B1 => inputs(73), B2 
                           => n15, ZN => n32);
   U43 : NAND4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => 
                           N133);
   U44 : AOI22_X1 port map( A1 => inputs(6), A2 => n10, B1 => inputs(108), B2 
                           => n3, ZN => n39);
   U45 : AOI22_X1 port map( A1 => inputs(23), A2 => n5, B1 => inputs(57), B2 =>
                           n11, ZN => n38);
   U46 : AOI22_X1 port map( A1 => inputs(40), A2 => n12, B1 => inputs(91), B2 
                           => n13, ZN => n37);
   U47 : AOI22_X1 port map( A1 => inputs(125), A2 => n14, B1 => inputs(74), B2 
                           => n15, ZN => n36);
   U48 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           N132);
   U49 : AOI22_X1 port map( A1 => inputs(7), A2 => n10, B1 => inputs(109), B2 
                           => n3, ZN => n43);
   U50 : AOI22_X1 port map( A1 => inputs(24), A2 => n5, B1 => inputs(58), B2 =>
                           n11, ZN => n42);
   U51 : AOI22_X1 port map( A1 => inputs(41), A2 => n12, B1 => inputs(92), B2 
                           => n13, ZN => n41);
   U52 : AOI22_X1 port map( A1 => inputs(126), A2 => n14, B1 => inputs(75), B2 
                           => n15, ZN => n40);
   U53 : NAND4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => 
                           N131);
   U54 : AOI22_X1 port map( A1 => inputs(8), A2 => n10, B1 => inputs(110), B2 
                           => n3, ZN => n47);
   U55 : AOI22_X1 port map( A1 => inputs(25), A2 => n5, B1 => inputs(59), B2 =>
                           n11, ZN => n46);
   U56 : AOI22_X1 port map( A1 => inputs(42), A2 => n12, B1 => inputs(93), B2 
                           => n13, ZN => n45);
   U57 : AOI22_X1 port map( A1 => inputs(127), A2 => n14, B1 => inputs(76), B2 
                           => n15, ZN => n44);
   U58 : NAND4_X1 port map( A1 => n48, A2 => n49, A3 => n50, A4 => n51, ZN => 
                           N130);
   U59 : AOI22_X1 port map( A1 => inputs(9), A2 => n10, B1 => inputs(111), B2 
                           => n3, ZN => n51);
   U60 : AOI22_X1 port map( A1 => inputs(26), A2 => n5, B1 => inputs(60), B2 =>
                           n11, ZN => n50);
   U61 : AOI22_X1 port map( A1 => inputs(43), A2 => n12, B1 => inputs(94), B2 
                           => n13, ZN => n49);
   U62 : AOI22_X1 port map( A1 => inputs(128), A2 => n14, B1 => inputs(77), B2 
                           => n15, ZN => n48);
   U63 : NAND4_X1 port map( A1 => n52, A2 => n53, A3 => n54, A4 => n55, ZN => 
                           N129);
   U64 : AOI22_X1 port map( A1 => inputs(10), A2 => n10, B1 => inputs(112), B2 
                           => n3, ZN => n55);
   U65 : AOI22_X1 port map( A1 => inputs(27), A2 => n5, B1 => inputs(61), B2 =>
                           n11, ZN => n54);
   U66 : AOI22_X1 port map( A1 => inputs(44), A2 => n12, B1 => inputs(95), B2 
                           => n13, ZN => n53);
   U67 : AOI22_X1 port map( A1 => inputs(129), A2 => n14, B1 => inputs(78), B2 
                           => n15, ZN => n52);
   U68 : NAND4_X1 port map( A1 => n56, A2 => n57, A3 => n58, A4 => n59, ZN => 
                           N128);
   U69 : AOI22_X1 port map( A1 => inputs(11), A2 => n10, B1 => inputs(113), B2 
                           => n3, ZN => n59);
   U70 : AOI22_X1 port map( A1 => inputs(28), A2 => n5, B1 => inputs(62), B2 =>
                           n11, ZN => n58);
   U71 : AOI22_X1 port map( A1 => inputs(45), A2 => n12, B1 => inputs(96), B2 
                           => n13, ZN => n57);
   U72 : AOI22_X1 port map( A1 => inputs(130), A2 => n14, B1 => inputs(79), B2 
                           => n15, ZN => n56);
   U73 : NAND4_X1 port map( A1 => n60, A2 => n61, A3 => n62, A4 => n63, ZN => 
                           N127);
   U74 : AOI22_X1 port map( A1 => inputs(12), A2 => n10, B1 => inputs(114), B2 
                           => n3, ZN => n63);
   U75 : AOI22_X1 port map( A1 => inputs(29), A2 => n5, B1 => inputs(63), B2 =>
                           n11, ZN => n62);
   U76 : AOI22_X1 port map( A1 => inputs(46), A2 => n12, B1 => inputs(97), B2 
                           => n13, ZN => n61);
   U77 : AOI22_X1 port map( A1 => inputs(131), A2 => n14, B1 => inputs(80), B2 
                           => n15, ZN => n60);
   U78 : NAND4_X1 port map( A1 => n64, A2 => n65, A3 => n66, A4 => n67, ZN => 
                           N126);
   U79 : AOI22_X1 port map( A1 => inputs(13), A2 => n10, B1 => inputs(115), B2 
                           => n3, ZN => n67);
   U80 : AOI22_X1 port map( A1 => inputs(30), A2 => n5, B1 => inputs(64), B2 =>
                           n11, ZN => n66);
   U81 : AOI22_X1 port map( A1 => inputs(47), A2 => n12, B1 => inputs(98), B2 
                           => n13, ZN => n65);
   U82 : AOI22_X1 port map( A1 => inputs(132), A2 => n14, B1 => inputs(81), B2 
                           => n15, ZN => n64);
   U83 : NAND4_X1 port map( A1 => n68, A2 => n69, A3 => n70, A4 => n71, ZN => 
                           N125);
   U84 : AOI22_X1 port map( A1 => inputs(14), A2 => n10, B1 => inputs(116), B2 
                           => n3, ZN => n71);
   U85 : AOI22_X1 port map( A1 => inputs(31), A2 => n5, B1 => inputs(65), B2 =>
                           n11, ZN => n70);
   U86 : AOI22_X1 port map( A1 => inputs(48), A2 => n12, B1 => inputs(99), B2 
                           => n13, ZN => n69);
   U87 : AOI22_X1 port map( A1 => inputs(133), A2 => n14, B1 => inputs(82), B2 
                           => n15, ZN => n68);
   U88 : NAND4_X1 port map( A1 => n72, A2 => n73, A3 => n74, A4 => n75, ZN => 
                           N124);
   U89 : AOI22_X1 port map( A1 => inputs(15), A2 => n10, B1 => inputs(117), B2 
                           => n3, ZN => n75);
   U90 : AOI22_X1 port map( A1 => inputs(32), A2 => n5, B1 => inputs(66), B2 =>
                           n11, ZN => n74);
   U91 : AOI22_X1 port map( A1 => inputs(49), A2 => n12, B1 => inputs(100), B2 
                           => n13, ZN => n73);
   U92 : AOI22_X1 port map( A1 => inputs(134), A2 => n14, B1 => inputs(83), B2 
                           => n15, ZN => n72);
   U93 : NAND4_X1 port map( A1 => n76, A2 => n77, A3 => n78, A4 => n79, ZN => 
                           N123);
   U94 : AOI22_X1 port map( A1 => inputs(16), A2 => n10, B1 => inputs(118), B2 
                           => n3, ZN => n79);
   U95 : OR4_X1 port map( A1 => n15, A2 => n14, A3 => n13, A4 => n12, ZN => n80
                           );
   U96 : AOI22_X1 port map( A1 => inputs(33), A2 => n5, B1 => inputs(67), B2 =>
                           n11, ZN => n78);
   U97 : AOI22_X1 port map( A1 => inputs(50), A2 => n12, B1 => inputs(101), B2 
                           => n13, ZN => n77);
   U98 : AOI22_X1 port map( A1 => inputs(135), A2 => n14, B1 => inputs(84), B2 
                           => n15, ZN => n76);
   U99 : INV_X1 port map( A => SEL(1), ZN => n82);
   U101 : INV_X1 port map( A => SEL(2), ZN => n81);
   U102 : INV_X1 port map( A => SEL(0), ZN => n83);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity encoder_0 is

   port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end encoder_0;

architecture SYN_beh of encoder_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_2_port, sel_1_port, sel_0_port, n1, n2, n3 : std_logic;

begin
   sel <= ( sel_2_port, sel_1_port, sel_0_port );
   
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => sel_1_port);
   U4 : NAND3_X1 port map( A1 => y(0), A2 => n3, A3 => y(1), ZN => n2);
   U5 : INV_X1 port map( A => sel_2_port, ZN => n1);
   U6 : AOI21_X1 port map( B1 => y(0), B2 => y(1), A => n3, ZN => sel_2_port);
   U7 : INV_X1 port map( A => y(2), ZN => n3);
   U8 : XOR2_X1 port map( A => y(1), B => y(0), Z => sel_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity complement2_N17 is

   port( value_in : in std_logic_vector (16 downto 0);  value_out : out 
         std_logic_vector (16 downto 0));

end complement2_N17;

architecture SYN_beh of complement2_N17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complement2_N17_DW01_inc_0
      port( A : in std_logic_vector (16 downto 0);  SUM : out std_logic_vector 
            (16 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N16, N15, N14, N13, N12, N11, N10, N1
      , N0 : std_logic;

begin
   
   add_0_root_add_22_ni : complement2_N17_DW01_inc_0 port map( A(16) => N0, 
                           A(15) => N1, A(14) => N2, A(13) => N3, A(12) => N4, 
                           A(11) => N5, A(10) => N6, A(9) => N7, A(8) => N8, 
                           A(7) => N9, A(6) => N10, A(5) => N11, A(4) => N12, 
                           A(3) => N13, A(2) => N14, A(1) => N15, A(0) => N16, 
                           SUM(16) => value_out(16), SUM(15) => value_out(15), 
                           SUM(14) => value_out(14), SUM(13) => value_out(13), 
                           SUM(12) => value_out(12), SUM(11) => value_out(11), 
                           SUM(10) => value_out(10), SUM(9) => value_out(9), 
                           SUM(8) => value_out(8), SUM(7) => value_out(7), 
                           SUM(6) => value_out(6), SUM(5) => value_out(5), 
                           SUM(4) => value_out(4), SUM(3) => value_out(3), 
                           SUM(2) => value_out(2), SUM(1) => value_out(1), 
                           SUM(0) => value_out(0));
   U2 : INV_X1 port map( A => value_in(7), ZN => N9);
   U3 : INV_X1 port map( A => value_in(8), ZN => N8);
   U4 : INV_X1 port map( A => value_in(9), ZN => N7);
   U5 : INV_X1 port map( A => value_in(10), ZN => N6);
   U6 : INV_X1 port map( A => value_in(11), ZN => N5);
   U7 : INV_X1 port map( A => value_in(12), ZN => N4);
   U8 : INV_X1 port map( A => value_in(13), ZN => N3);
   U9 : INV_X1 port map( A => value_in(14), ZN => N2);
   U10 : INV_X1 port map( A => value_in(0), ZN => N16);
   U11 : INV_X1 port map( A => value_in(1), ZN => N15);
   U12 : INV_X1 port map( A => value_in(2), ZN => N14);
   U13 : INV_X1 port map( A => value_in(3), ZN => N13);
   U14 : INV_X1 port map( A => value_in(4), ZN => N12);
   U15 : INV_X1 port map( A => value_in(5), ZN => N11);
   U16 : INV_X1 port map( A => value_in(6), ZN => N10);
   U17 : INV_X1 port map( A => value_in(15), ZN => N1);
   U18 : INV_X1 port map( A => value_in(16), ZN => N0);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SUM_GEN_NBIT32_NBLOCKS4 is

   port( A, B, Ci : in std_logic_vector (31 downto 0);  S : out 
         std_logic_vector (31 downto 0));

end SUM_GEN_NBIT32_NBLOCKS4;

architecture SYN_STRUCTURAL of SUM_GEN_NBIT32_NBLOCKS4 is

   component CSB_NBIT8_1
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component CSB_NBIT8_2
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component CSB_NBIT8_3
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component CSB_NBIT8_0
      port( A, B : in std_logic_vector (7 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (7 downto 0));
   end component;

begin
   
   CSBi_0 : CSB_NBIT8_0 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(7) => B(7), B(6) => B(6), B(5)
                           => B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), Ci => Ci(0), S(7) => 
                           S(7), S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3)
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBi_1 : CSB_NBIT8_3 port map( A(7) => A(15), A(6) => A(14), A(5) => A(13), 
                           A(4) => A(12), A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(7) => B(15), B(6) => B(14), 
                           B(5) => B(13), B(4) => B(12), B(3) => B(11), B(2) =>
                           B(10), B(1) => B(9), B(0) => B(8), Ci => Ci(8), S(7)
                           => S(15), S(6) => S(14), S(5) => S(13), S(4) => 
                           S(12), S(3) => S(11), S(2) => S(10), S(1) => S(9), 
                           S(0) => S(8));
   CSBi_2 : CSB_NBIT8_2 port map( A(7) => A(23), A(6) => A(22), A(5) => A(21), 
                           A(4) => A(20), A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(7) => B(23), B(6) => B(22), 
                           B(5) => B(21), B(4) => B(20), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Ci(16), 
                           S(7) => S(23), S(6) => S(22), S(5) => S(21), S(4) =>
                           S(20), S(3) => S(19), S(2) => S(18), S(1) => S(17), 
                           S(0) => S(16));
   CSBi_3 : CSB_NBIT8_1 port map( A(7) => A(31), A(6) => A(30), A(5) => A(29), 
                           A(4) => A(28), A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(7) => B(31), B(6) => B(30), 
                           B(5) => B(29), B(4) => B(28), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Ci(24), 
                           S(7) => S(31), S(6) => S(30), S(5) => S(29), S(4) =>
                           S(28), S(3) => S(27), S(2) => S(26), S(1) => S(25), 
                           S(0) => S(24));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity STCG_NBIT32_SDIST4 is

   port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  Cout :
         out std_logic_vector (32 downto 0));

end STCG_NBIT32_SDIST4;

architecture SYN_STRUCTURAL of STCG_NBIT32_SDIST4 is

   component GSB_1
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component GSB_2
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component GSB_3
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component GSB_4
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component PGSB_1
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_2
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GSB_5
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component GSB_6
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component PGSB_3
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_4
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_5
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GSB_7
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component PGSB_6
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_7
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_8
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_9
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_10
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_11
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_12
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GSB_8
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component PGSB_13
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_14
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_15
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_16
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_17
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_18
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_19
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_20
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_21
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_22
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_23
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_24
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_25
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_26
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component PGSB_0
      port( P_in_ik, P_in_kj, G_in_ik, G_in_kj : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GSB_0
      port( P_in_ik, G_in_ik, G_in_kj : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  p, 
            g : out std_logic_vector (31 downto 0));
   end component;
   
   signal Cout_32_port, Cout_28, Cout_24, Cout_20, Cout_16, Cout_12, Cout_8, 
      Cout_4, g_4_31_port, g_4_27_port, g_3_31_port, g_3_23_port, g_3_15_port, 
      g_2_31_port, g_2_27_port, g_2_23_port, g_2_19_port, g_2_15_port, 
      g_2_11_port, g_2_7_port, g_1_31_port, g_1_29_port, g_1_27_port, 
      g_1_25_port, g_1_23_port, g_1_21_port, g_1_19_port, g_1_17_port, 
      g_1_15_port, g_1_13_port, g_1_11_port, g_1_9_port, g_1_7_port, g_1_5_port
      , g_1_3_port, g_1_1_port, g_0_31_port, g_0_30_port, g_0_29_port, 
      g_0_28_port, g_0_27_port, g_0_26_port, g_0_25_port, g_0_24_port, 
      g_0_23_port, g_0_22_port, g_0_21_port, g_0_20_port, g_0_19_port, 
      g_0_18_port, g_0_17_port, g_0_16_port, g_0_15_port, g_0_14_port, 
      g_0_13_port, g_0_12_port, g_0_11_port, g_0_10_port, g_0_9_port, 
      g_0_8_port, g_0_7_port, g_0_6_port, g_0_5_port, g_0_4_port, g_0_3_port, 
      g_0_2_port, g_0_1_port, g_0_0_port, p_4_31_port, p_4_27_port, p_3_31_port
      , p_3_23_port, p_3_15_port, p_2_31_port, p_2_27_port, p_2_23_port, 
      p_2_19_port, p_2_15_port, p_2_11_port, p_2_7_port, p_1_31_port, 
      p_1_29_port, p_1_27_port, p_1_25_port, p_1_23_port, p_1_21_port, 
      p_1_19_port, p_1_17_port, p_1_15_port, p_1_13_port, p_1_11_port, 
      p_1_9_port, p_1_7_port, p_1_5_port, p_1_3_port, p_0_31_port, p_0_30_port,
      p_0_29_port, p_0_28_port, p_0_27_port, p_0_26_port, p_0_25_port, 
      p_0_24_port, p_0_23_port, p_0_22_port, p_0_21_port, p_0_20_port, 
      p_0_19_port, p_0_18_port, p_0_17_port, p_0_16_port, p_0_15_port, 
      p_0_14_port, p_0_13_port, p_0_12_port, p_0_11_port, p_0_10_port, 
      p_0_9_port, p_0_8_port, p_0_7_port, p_0_6_port, p_0_5_port, p_0_4_port, 
      p_0_3_port, p_0_2_port, p_0_1_port, net5404, net5405, net5406, net5407, 
      net5408, net5409, net5410, net5411, net5412, net5413, net5414, net5415, 
      net5416, net5417, net5418, net5419, net5420, net5421, net5422, net5423, 
      net5424, net5425, net5426, net5427, n_3356 : std_logic;

begin
   Cout <= ( Cout_32_port, net5427, net5426, net5425, Cout_28, net5424, net5423
      , net5422, Cout_24, net5421, net5420, net5419, Cout_20, net5418, net5417,
      net5416, Cout_16, net5415, net5414, net5413, Cout_12, net5412, net5411, 
      net5410, Cout_8, net5409, net5408, net5407, Cout_4, net5406, net5405, 
      net5404, cin );
   
   net5404 <= '0';
   net5405 <= '0';
   net5406 <= '0';
   net5407 <= '0';
   net5408 <= '0';
   net5409 <= '0';
   net5410 <= '0';
   net5411 <= '0';
   net5412 <= '0';
   net5413 <= '0';
   net5414 <= '0';
   net5415 <= '0';
   net5416 <= '0';
   net5417 <= '0';
   net5418 <= '0';
   net5419 <= '0';
   net5420 <= '0';
   net5421 <= '0';
   net5422 <= '0';
   net5423 <= '0';
   net5424 <= '0';
   net5425 <= '0';
   net5426 <= '0';
   net5427 <= '0';
   PGnetwork : PG_NBIT32 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), cin => cin, p(31) => p_0_31_port, p(30) => 
                           p_0_30_port, p(29) => p_0_29_port, p(28) => 
                           p_0_28_port, p(27) => p_0_27_port, p(26) => 
                           p_0_26_port, p(25) => p_0_25_port, p(24) => 
                           p_0_24_port, p(23) => p_0_23_port, p(22) => 
                           p_0_22_port, p(21) => p_0_21_port, p(20) => 
                           p_0_20_port, p(19) => p_0_19_port, p(18) => 
                           p_0_18_port, p(17) => p_0_17_port, p(16) => 
                           p_0_16_port, p(15) => p_0_15_port, p(14) => 
                           p_0_14_port, p(13) => p_0_13_port, p(12) => 
                           p_0_12_port, p(11) => p_0_11_port, p(10) => 
                           p_0_10_port, p(9) => p_0_9_port, p(8) => p_0_8_port,
                           p(7) => p_0_7_port, p(6) => p_0_6_port, p(5) => 
                           p_0_5_port, p(4) => p_0_4_port, p(3) => p_0_3_port, 
                           p(2) => p_0_2_port, p(1) => p_0_1_port, p(0) => 
                           n_3356, g(31) => g_0_31_port, g(30) => g_0_30_port, 
                           g(29) => g_0_29_port, g(28) => g_0_28_port, g(27) =>
                           g_0_27_port, g(26) => g_0_26_port, g(25) => 
                           g_0_25_port, g(24) => g_0_24_port, g(23) => 
                           g_0_23_port, g(22) => g_0_22_port, g(21) => 
                           g_0_21_port, g(20) => g_0_20_port, g(19) => 
                           g_0_19_port, g(18) => g_0_18_port, g(17) => 
                           g_0_17_port, g(16) => g_0_16_port, g(15) => 
                           g_0_15_port, g(14) => g_0_14_port, g(13) => 
                           g_0_13_port, g(12) => g_0_12_port, g(11) => 
                           g_0_11_port, g(10) => g_0_10_port, g(9) => 
                           g_0_9_port, g(8) => g_0_8_port, g(7) => g_0_7_port, 
                           g(6) => g_0_6_port, g(5) => g_0_5_port, g(4) => 
                           g_0_4_port, g(3) => g_0_3_port, g(2) => g_0_2_port, 
                           g(1) => g_0_1_port, g(0) => g_0_0_port);
   Gi_1_1 : GSB_0 port map( P_in_ik => p_0_1_port, G_in_ik => g_0_1_port, 
                           G_in_kj => g_0_0_port, G_out => g_1_1_port);
   PGi_1_3 : PGSB_0 port map( P_in_ik => p_0_3_port, P_in_kj => p_0_2_port, 
                           G_in_ik => g_0_3_port, G_in_kj => g_0_2_port, G_out 
                           => g_1_3_port, P_out => p_1_3_port);
   PGi_1_5 : PGSB_26 port map( P_in_ik => p_0_5_port, P_in_kj => p_0_4_port, 
                           G_in_ik => g_0_5_port, G_in_kj => g_0_4_port, G_out 
                           => g_1_5_port, P_out => p_1_5_port);
   PGi_1_7 : PGSB_25 port map( P_in_ik => p_0_7_port, P_in_kj => p_0_6_port, 
                           G_in_ik => g_0_7_port, G_in_kj => g_0_6_port, G_out 
                           => g_1_7_port, P_out => p_1_7_port);
   PGi_1_9 : PGSB_24 port map( P_in_ik => p_0_9_port, P_in_kj => p_0_8_port, 
                           G_in_ik => g_0_9_port, G_in_kj => g_0_8_port, G_out 
                           => g_1_9_port, P_out => p_1_9_port);
   PGi_1_11 : PGSB_23 port map( P_in_ik => p_0_11_port, P_in_kj => p_0_10_port,
                           G_in_ik => g_0_11_port, G_in_kj => g_0_10_port, 
                           G_out => g_1_11_port, P_out => p_1_11_port);
   PGi_1_13 : PGSB_22 port map( P_in_ik => p_0_13_port, P_in_kj => p_0_12_port,
                           G_in_ik => g_0_13_port, G_in_kj => g_0_12_port, 
                           G_out => g_1_13_port, P_out => p_1_13_port);
   PGi_1_15 : PGSB_21 port map( P_in_ik => p_0_15_port, P_in_kj => p_0_14_port,
                           G_in_ik => g_0_15_port, G_in_kj => g_0_14_port, 
                           G_out => g_1_15_port, P_out => p_1_15_port);
   PGi_1_17 : PGSB_20 port map( P_in_ik => p_0_17_port, P_in_kj => p_0_16_port,
                           G_in_ik => g_0_17_port, G_in_kj => g_0_16_port, 
                           G_out => g_1_17_port, P_out => p_1_17_port);
   PGi_1_19 : PGSB_19 port map( P_in_ik => p_0_19_port, P_in_kj => p_0_18_port,
                           G_in_ik => g_0_19_port, G_in_kj => g_0_18_port, 
                           G_out => g_1_19_port, P_out => p_1_19_port);
   PGi_1_21 : PGSB_18 port map( P_in_ik => p_0_21_port, P_in_kj => p_0_20_port,
                           G_in_ik => g_0_21_port, G_in_kj => g_0_20_port, 
                           G_out => g_1_21_port, P_out => p_1_21_port);
   PGi_1_23 : PGSB_17 port map( P_in_ik => p_0_23_port, P_in_kj => p_0_22_port,
                           G_in_ik => g_0_23_port, G_in_kj => g_0_22_port, 
                           G_out => g_1_23_port, P_out => p_1_23_port);
   PGi_1_25 : PGSB_16 port map( P_in_ik => p_0_25_port, P_in_kj => p_0_24_port,
                           G_in_ik => g_0_25_port, G_in_kj => g_0_24_port, 
                           G_out => g_1_25_port, P_out => p_1_25_port);
   PGi_1_27 : PGSB_15 port map( P_in_ik => p_0_27_port, P_in_kj => p_0_26_port,
                           G_in_ik => g_0_27_port, G_in_kj => g_0_26_port, 
                           G_out => g_1_27_port, P_out => p_1_27_port);
   PGi_1_29 : PGSB_14 port map( P_in_ik => p_0_29_port, P_in_kj => p_0_28_port,
                           G_in_ik => g_0_29_port, G_in_kj => g_0_28_port, 
                           G_out => g_1_29_port, P_out => p_1_29_port);
   PGi_1_31 : PGSB_13 port map( P_in_ik => p_0_31_port, P_in_kj => p_0_30_port,
                           G_in_ik => g_0_31_port, G_in_kj => g_0_30_port, 
                           G_out => g_1_31_port, P_out => p_1_31_port);
   Gi_2_3 : GSB_8 port map( P_in_ik => p_1_3_port, G_in_ik => g_1_3_port, 
                           G_in_kj => g_1_1_port, G_out => Cout_4);
   PGi_2_7 : PGSB_12 port map( P_in_ik => p_1_7_port, P_in_kj => p_1_5_port, 
                           G_in_ik => g_1_7_port, G_in_kj => g_1_5_port, G_out 
                           => g_2_7_port, P_out => p_2_7_port);
   PGi_2_11 : PGSB_11 port map( P_in_ik => p_1_11_port, P_in_kj => p_1_9_port, 
                           G_in_ik => g_1_11_port, G_in_kj => g_1_9_port, G_out
                           => g_2_11_port, P_out => p_2_11_port);
   PGi_2_15 : PGSB_10 port map( P_in_ik => p_1_15_port, P_in_kj => p_1_13_port,
                           G_in_ik => g_1_15_port, G_in_kj => g_1_13_port, 
                           G_out => g_2_15_port, P_out => p_2_15_port);
   PGi_2_19 : PGSB_9 port map( P_in_ik => p_1_19_port, P_in_kj => p_1_17_port, 
                           G_in_ik => g_1_19_port, G_in_kj => g_1_17_port, 
                           G_out => g_2_19_port, P_out => p_2_19_port);
   PGi_2_23 : PGSB_8 port map( P_in_ik => p_1_23_port, P_in_kj => p_1_21_port, 
                           G_in_ik => g_1_23_port, G_in_kj => g_1_21_port, 
                           G_out => g_2_23_port, P_out => p_2_23_port);
   PGi_2_27 : PGSB_7 port map( P_in_ik => p_1_27_port, P_in_kj => p_1_25_port, 
                           G_in_ik => g_1_27_port, G_in_kj => g_1_25_port, 
                           G_out => g_2_27_port, P_out => p_2_27_port);
   PGi_2_31 : PGSB_6 port map( P_in_ik => p_1_31_port, P_in_kj => p_1_29_port, 
                           G_in_ik => g_1_31_port, G_in_kj => g_1_29_port, 
                           G_out => g_2_31_port, P_out => p_2_31_port);
   Gi_3_7 : GSB_7 port map( P_in_ik => p_2_7_port, G_in_ik => g_2_7_port, 
                           G_in_kj => Cout_4, G_out => Cout_8);
   PGi_3_15 : PGSB_5 port map( P_in_ik => p_2_15_port, P_in_kj => p_2_11_port, 
                           G_in_ik => g_2_15_port, G_in_kj => g_2_11_port, 
                           G_out => g_3_15_port, P_out => p_3_15_port);
   PGi_3_23 : PGSB_4 port map( P_in_ik => p_2_23_port, P_in_kj => p_2_19_port, 
                           G_in_ik => g_2_23_port, G_in_kj => g_2_19_port, 
                           G_out => g_3_23_port, P_out => p_3_23_port);
   PGi_3_31 : PGSB_3 port map( P_in_ik => p_2_31_port, P_in_kj => p_2_27_port, 
                           G_in_ik => g_2_31_port, G_in_kj => g_2_27_port, 
                           G_out => g_3_31_port, P_out => p_3_31_port);
   Gi_4_11 : GSB_6 port map( P_in_ik => p_2_11_port, G_in_ik => g_2_11_port, 
                           G_in_kj => Cout_8, G_out => Cout_12);
   Gi_4_15 : GSB_5 port map( P_in_ik => p_3_15_port, G_in_ik => g_3_15_port, 
                           G_in_kj => Cout_8, G_out => Cout_16);
   PGi_4_27 : PGSB_2 port map( P_in_ik => p_2_27_port, P_in_kj => p_3_23_port, 
                           G_in_ik => g_2_27_port, G_in_kj => g_3_23_port, 
                           G_out => g_4_27_port, P_out => p_4_27_port);
   PGi_4_31 : PGSB_1 port map( P_in_ik => p_3_31_port, P_in_kj => p_3_23_port, 
                           G_in_ik => g_3_31_port, G_in_kj => g_3_23_port, 
                           G_out => g_4_31_port, P_out => p_4_31_port);
   Gi_5_19 : GSB_4 port map( P_in_ik => p_2_19_port, G_in_ik => g_2_19_port, 
                           G_in_kj => Cout_16, G_out => Cout_20);
   Gi_5_23 : GSB_3 port map( P_in_ik => p_3_23_port, G_in_ik => g_3_23_port, 
                           G_in_kj => Cout_16, G_out => Cout_24);
   Gi_5_27 : GSB_2 port map( P_in_ik => p_4_27_port, G_in_ik => g_4_27_port, 
                           G_in_kj => Cout_16, G_out => Cout_28);
   Gi_5_31 : GSB_1 port map( P_in_ik => p_4_31_port, G_in_ik => g_4_31_port, 
                           G_in_kj => Cout_16, G_out => Cout_32_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity boothmul_pipelined_N16 is

   port( clk, rst : in std_logic;  multiplier, multiplicand : in 
         std_logic_vector (15 downto 0);  result : out std_logic_vector (31 
         downto 0));

end boothmul_pipelined_N16;

architecture SYN_struc of boothmul_pipelined_N16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component reg_nbit_n16_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component reg_nbit_n16_2
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component reg_nbit_n16_3
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component reg_nbit_n16_4
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component reg_nbit_n16_5
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component reg_nbit_n16_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (15 downto 0); 
            Q : out std_logic_vector (15 downto 0));
   end component;
   
   component adder_NBIT31
      port( a, b : in std_logic_vector (30 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX_zbit_nbit_N31_Z3
      port( inputs : in std_logic_vector (0 to 247);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (30 downto 0));
   end component;
   
   component reg_nbit_n249_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_1
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT29
      port( a, b : in std_logic_vector (28 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (29 downto 0));
   end component;
   
   component MUX_zbit_nbit_N29_Z3
      port( inputs : in std_logic_vector (0 to 231);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (28 downto 0));
   end component;
   
   component reg_nbit_n249_2
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_2
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_2
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT27
      port( a, b : in std_logic_vector (26 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (27 downto 0));
   end component;
   
   component MUX_zbit_nbit_N27_Z3
      port( inputs : in std_logic_vector (0 to 215);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (26 downto 0));
   end component;
   
   component reg_nbit_n249_3
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_3
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_3
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT25
      port( a, b : in std_logic_vector (24 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (25 downto 0));
   end component;
   
   component MUX_zbit_nbit_N25_Z3
      port( inputs : in std_logic_vector (0 to 199);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (24 downto 0));
   end component;
   
   component reg_nbit_n249_4
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_4
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_4
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT23
      port( a, b : in std_logic_vector (22 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (23 downto 0));
   end component;
   
   component MUX_zbit_nbit_N23_Z3
      port( inputs : in std_logic_vector (0 to 183);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (22 downto 0));
   end component;
   
   component reg_nbit_n249_5
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_5
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_5
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT21
      port( a, b : in std_logic_vector (20 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (21 downto 0));
   end component;
   
   component MUX_zbit_nbit_N21_Z3
      port( inputs : in std_logic_vector (0 to 167);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (20 downto 0));
   end component;
   
   component reg_nbit_n249_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (248 downto 0);
            Q : out std_logic_vector (248 downto 0));
   end component;
   
   component encoder_6
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component reg_nbit_n32_6
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT19
      port( a, b : in std_logic_vector (18 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (19 downto 0));
   end component;
   
   component MUX_zbit_nbit_N19_Z3
      port( inputs : in std_logic_vector (0 to 151);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (18 downto 0));
   end component;
   
   component encoder_7
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_zbit_nbit_N17_Z3
      port( inputs : in std_logic_vector (0 to 135);  SEL : in std_logic_vector
            (2 downto 0);  Y : out std_logic_vector (16 downto 0));
   end component;
   
   component encoder_0
      port( y : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component complement2_N17
      port( value_in : in std_logic_vector (16 downto 0);  value_out : out 
            std_logic_vector (16 downto 0));
   end component;
   
   signal X_Logic0_port, muxes_in_0_102_port, muxes_in_0_103_port, 
      muxes_in_0_104_port, muxes_in_0_105_port, muxes_in_0_106_port, 
      muxes_in_0_107_port, muxes_in_0_108_port, muxes_in_0_109_port, 
      muxes_in_0_110_port, muxes_in_0_111_port, muxes_in_0_112_port, 
      muxes_in_0_113_port, muxes_in_0_114_port, muxes_in_0_115_port, 
      muxes_in_0_116_port, muxes_in_0_117_port, muxes_in_0_119_port, 
      multiplicand_pip_2_15_port, multiplicand_pip_2_14_port, 
      multiplicand_pip_2_13_port, multiplicand_pip_2_12_port, 
      multiplicand_pip_2_11_port, multiplicand_pip_2_10_port, 
      multiplicand_pip_2_9_port, multiplicand_pip_2_8_port, 
      multiplicand_pip_2_7_port, multiplicand_pip_2_6_port, 
      multiplicand_pip_2_5_port, multiplicand_pip_2_4_port, 
      multiplicand_pip_2_3_port, multiplicand_pip_2_2_port, 
      multiplicand_pip_2_1_port, multiplicand_pip_2_0_port, 
      multiplicand_pip_3_15_port, multiplicand_pip_3_14_port, 
      multiplicand_pip_3_13_port, multiplicand_pip_3_12_port, 
      multiplicand_pip_3_11_port, multiplicand_pip_3_10_port, 
      multiplicand_pip_3_9_port, multiplicand_pip_3_8_port, 
      multiplicand_pip_3_7_port, multiplicand_pip_3_6_port, 
      multiplicand_pip_3_5_port, multiplicand_pip_3_4_port, 
      multiplicand_pip_3_3_port, multiplicand_pip_3_2_port, 
      multiplicand_pip_3_1_port, multiplicand_pip_3_0_port, 
      multiplicand_pip_4_15_port, multiplicand_pip_4_14_port, 
      multiplicand_pip_4_13_port, multiplicand_pip_4_12_port, 
      multiplicand_pip_4_11_port, multiplicand_pip_4_10_port, 
      multiplicand_pip_4_9_port, multiplicand_pip_4_8_port, 
      multiplicand_pip_4_7_port, multiplicand_pip_4_6_port, 
      multiplicand_pip_4_5_port, multiplicand_pip_4_4_port, 
      multiplicand_pip_4_3_port, multiplicand_pip_4_2_port, 
      multiplicand_pip_4_1_port, multiplicand_pip_4_0_port, 
      multiplicand_pip_5_15_port, multiplicand_pip_5_14_port, 
      multiplicand_pip_5_13_port, multiplicand_pip_5_12_port, 
      multiplicand_pip_5_11_port, multiplicand_pip_5_10_port, 
      multiplicand_pip_5_9_port, multiplicand_pip_5_8_port, 
      multiplicand_pip_5_7_port, multiplicand_pip_5_6_port, 
      multiplicand_pip_5_5_port, multiplicand_pip_5_4_port, 
      multiplicand_pip_5_3_port, multiplicand_pip_5_2_port, 
      multiplicand_pip_5_1_port, multiplicand_pip_5_0_port, 
      multiplicand_pip_6_15_port, multiplicand_pip_6_14_port, 
      multiplicand_pip_6_13_port, multiplicand_pip_6_12_port, 
      multiplicand_pip_6_11_port, multiplicand_pip_6_10_port, 
      multiplicand_pip_6_9_port, multiplicand_pip_6_8_port, 
      multiplicand_pip_6_7_port, multiplicand_pip_6_6_port, 
      multiplicand_pip_6_5_port, multiplicand_pip_6_4_port, 
      multiplicand_pip_6_3_port, multiplicand_pip_6_2_port, 
      multiplicand_pip_6_1_port, multiplicand_pip_6_0_port, 
      multiplicand_pip_7_15_port, multiplicand_pip_7_14_port, 
      multiplicand_pip_7_13_port, encoder_out_0_2_port, encoder_out_0_1_port, 
      encoder_out_0_0_port, encoder_out_1_2_port, encoder_out_1_1_port, 
      encoder_out_1_0_port, encoder_out_2_2_port, encoder_out_2_1_port, 
      encoder_out_2_0_port, encoder_out_3_2_port, encoder_out_3_1_port, 
      encoder_out_3_0_port, encoder_out_4_2_port, encoder_out_4_1_port, 
      encoder_out_4_0_port, encoder_out_5_2_port, encoder_out_5_1_port, 
      encoder_out_5_0_port, encoder_out_6_2_port, encoder_out_6_1_port, 
      encoder_out_6_0_port, encoder_out_7_2_port, encoder_out_7_1_port, 
      encoder_out_7_0_port, mux_out_1_18_port, mux_out_1_17_port, 
      mux_out_1_16_port, mux_out_1_15_port, mux_out_1_14_port, 
      mux_out_1_13_port, mux_out_1_12_port, mux_out_1_11_port, 
      mux_out_1_10_port, mux_out_1_9_port, mux_out_1_8_port, mux_out_1_7_port, 
      mux_out_1_6_port, mux_out_1_5_port, mux_out_1_4_port, mux_out_1_3_port, 
      mux_out_1_2_port, mux_out_1_1_port, mux_out_1_0_port, mux_out_2_20_port, 
      mux_out_2_19_port, mux_out_2_18_port, mux_out_2_17_port, 
      mux_out_2_16_port, mux_out_2_15_port, mux_out_2_14_port, 
      mux_out_2_13_port, mux_out_2_12_port, mux_out_2_11_port, 
      mux_out_2_10_port, mux_out_2_9_port, mux_out_2_8_port, mux_out_2_7_port, 
      mux_out_2_6_port, mux_out_2_5_port, mux_out_2_4_port, mux_out_2_3_port, 
      mux_out_2_2_port, mux_out_2_1_port, mux_out_2_0_port, mux_out_3_22_port, 
      mux_out_3_21_port, mux_out_3_20_port, mux_out_3_19_port, 
      mux_out_3_18_port, mux_out_3_17_port, mux_out_3_16_port, 
      mux_out_3_15_port, mux_out_3_14_port, mux_out_3_13_port, 
      mux_out_3_12_port, mux_out_3_11_port, mux_out_3_10_port, mux_out_3_9_port
      , mux_out_3_8_port, mux_out_3_7_port, mux_out_3_6_port, mux_out_3_5_port,
      mux_out_3_4_port, mux_out_3_3_port, mux_out_3_2_port, mux_out_3_1_port, 
      mux_out_3_0_port, mux_out_4_24_port, mux_out_4_23_port, mux_out_4_22_port
      , mux_out_4_21_port, mux_out_4_20_port, mux_out_4_19_port, 
      mux_out_4_18_port, mux_out_4_17_port, mux_out_4_16_port, 
      mux_out_4_15_port, mux_out_4_14_port, mux_out_4_13_port, 
      mux_out_4_12_port, mux_out_4_11_port, mux_out_4_10_port, mux_out_4_9_port
      , mux_out_4_8_port, mux_out_4_7_port, mux_out_4_6_port, mux_out_4_5_port,
      mux_out_4_4_port, mux_out_4_3_port, mux_out_4_2_port, mux_out_4_1_port, 
      mux_out_4_0_port, mux_out_5_26_port, mux_out_5_25_port, mux_out_5_24_port
      , mux_out_5_23_port, mux_out_5_22_port, mux_out_5_21_port, 
      mux_out_5_20_port, mux_out_5_19_port, mux_out_5_18_port, 
      mux_out_5_17_port, mux_out_5_16_port, mux_out_5_15_port, 
      mux_out_5_14_port, mux_out_5_13_port, mux_out_5_12_port, 
      mux_out_5_11_port, mux_out_5_10_port, mux_out_5_9_port, mux_out_5_8_port,
      mux_out_5_7_port, mux_out_5_6_port, mux_out_5_5_port, mux_out_5_4_port, 
      mux_out_5_3_port, mux_out_5_2_port, mux_out_5_1_port, mux_out_5_0_port, 
      mux_out_6_28_port, mux_out_6_27_port, mux_out_6_26_port, 
      mux_out_6_25_port, mux_out_6_24_port, mux_out_6_23_port, 
      mux_out_6_22_port, mux_out_6_21_port, mux_out_6_20_port, 
      mux_out_6_19_port, mux_out_6_18_port, mux_out_6_17_port, 
      mux_out_6_16_port, mux_out_6_15_port, mux_out_6_14_port, 
      mux_out_6_13_port, mux_out_6_12_port, mux_out_6_11_port, 
      mux_out_6_10_port, mux_out_6_9_port, mux_out_6_8_port, mux_out_6_7_port, 
      mux_out_6_6_port, mux_out_6_5_port, mux_out_6_4_port, mux_out_6_3_port, 
      mux_out_6_2_port, mux_out_6_1_port, mux_out_6_0_port, mux_out_7_30_port, 
      mux_out_7_29_port, mux_out_7_28_port, mux_out_7_27_port, 
      mux_out_7_26_port, mux_out_7_25_port, mux_out_7_24_port, 
      mux_out_7_23_port, mux_out_7_22_port, mux_out_7_21_port, 
      mux_out_7_20_port, mux_out_7_19_port, mux_out_7_18_port, 
      mux_out_7_17_port, mux_out_7_16_port, mux_out_7_15_port, 
      mux_out_7_14_port, mux_out_7_13_port, mux_out_7_12_port, 
      mux_out_7_11_port, mux_out_7_10_port, mux_out_7_9_port, mux_out_7_8_port,
      mux_out_7_7_port, mux_out_7_6_port, mux_out_7_5_port, mux_out_7_4_port, 
      mux_out_7_3_port, mux_out_7_2_port, mux_out_7_1_port, mux_out_7_0_port, 
      sum_B_in_1_18_port, sum_B_in_1_15_port, sum_B_in_1_14_port, 
      sum_B_in_1_13_port, sum_B_in_1_12_port, sum_B_in_1_11_port, 
      sum_B_in_1_10_port, sum_B_in_1_9_port, sum_B_in_1_8_port, 
      sum_B_in_1_7_port, sum_B_in_1_6_port, sum_B_in_1_5_port, 
      sum_B_in_1_4_port, sum_B_in_1_3_port, sum_B_in_1_2_port, 
      sum_B_in_1_1_port, sum_B_in_1_0_port, sum_B_in_2_20_port, 
      sum_B_in_2_17_port, sum_B_in_2_16_port, sum_B_in_2_15_port, 
      sum_B_in_2_14_port, sum_B_in_2_13_port, sum_B_in_2_12_port, 
      sum_B_in_2_11_port, sum_B_in_2_10_port, sum_B_in_2_9_port, 
      sum_B_in_2_8_port, sum_B_in_2_7_port, sum_B_in_2_6_port, 
      sum_B_in_2_5_port, sum_B_in_2_4_port, sum_B_in_2_3_port, 
      sum_B_in_2_2_port, sum_B_in_2_1_port, sum_B_in_2_0_port, 
      sum_B_in_3_22_port, sum_B_in_3_19_port, sum_B_in_3_18_port, 
      sum_B_in_3_17_port, sum_B_in_3_16_port, sum_B_in_3_15_port, 
      sum_B_in_3_14_port, sum_B_in_3_13_port, sum_B_in_3_12_port, 
      sum_B_in_3_11_port, sum_B_in_3_10_port, sum_B_in_3_9_port, 
      sum_B_in_3_8_port, sum_B_in_3_7_port, sum_B_in_3_6_port, 
      sum_B_in_3_5_port, sum_B_in_3_4_port, sum_B_in_3_3_port, 
      sum_B_in_3_2_port, sum_B_in_3_1_port, sum_B_in_3_0_port, 
      sum_B_in_4_24_port, sum_B_in_4_21_port, sum_B_in_4_20_port, 
      sum_B_in_4_19_port, sum_B_in_4_18_port, sum_B_in_4_17_port, 
      sum_B_in_4_16_port, sum_B_in_4_15_port, sum_B_in_4_14_port, 
      sum_B_in_4_13_port, sum_B_in_4_12_port, sum_B_in_4_11_port, 
      sum_B_in_4_10_port, sum_B_in_4_9_port, sum_B_in_4_8_port, 
      sum_B_in_4_7_port, sum_B_in_4_6_port, sum_B_in_4_5_port, 
      sum_B_in_4_4_port, sum_B_in_4_3_port, sum_B_in_4_2_port, 
      sum_B_in_4_1_port, sum_B_in_4_0_port, sum_B_in_5_26_port, 
      sum_B_in_5_23_port, sum_B_in_5_22_port, sum_B_in_5_21_port, 
      sum_B_in_5_20_port, sum_B_in_5_19_port, sum_B_in_5_18_port, 
      sum_B_in_5_17_port, sum_B_in_5_16_port, sum_B_in_5_15_port, 
      sum_B_in_5_14_port, sum_B_in_5_13_port, sum_B_in_5_12_port, 
      sum_B_in_5_11_port, sum_B_in_5_10_port, sum_B_in_5_9_port, 
      sum_B_in_5_8_port, sum_B_in_5_7_port, sum_B_in_5_6_port, 
      sum_B_in_5_5_port, sum_B_in_5_4_port, sum_B_in_5_3_port, 
      sum_B_in_5_2_port, sum_B_in_5_1_port, sum_B_in_5_0_port, 
      sum_B_in_6_28_port, sum_B_in_6_25_port, sum_B_in_6_24_port, 
      sum_B_in_6_23_port, sum_B_in_6_22_port, sum_B_in_6_21_port, 
      sum_B_in_6_20_port, sum_B_in_6_19_port, sum_B_in_6_18_port, 
      sum_B_in_6_17_port, sum_B_in_6_16_port, sum_B_in_6_15_port, 
      sum_B_in_6_14_port, sum_B_in_6_13_port, sum_B_in_6_12_port, 
      sum_B_in_6_11_port, sum_B_in_6_10_port, sum_B_in_6_9_port, 
      sum_B_in_6_8_port, sum_B_in_6_7_port, sum_B_in_6_6_port, 
      sum_B_in_6_5_port, sum_B_in_6_4_port, sum_B_in_6_3_port, 
      sum_B_in_6_2_port, sum_B_in_6_1_port, sum_B_in_6_0_port, 
      sum_B_in_7_30_port, sum_B_in_7_27_port, sum_B_in_7_26_port, 
      sum_B_in_7_25_port, sum_B_in_7_24_port, sum_B_in_7_23_port, 
      sum_B_in_7_22_port, sum_B_in_7_21_port, sum_B_in_7_20_port, 
      sum_B_in_7_19_port, sum_B_in_7_18_port, sum_B_in_7_17_port, 
      sum_B_in_7_16_port, sum_B_in_7_15_port, sum_B_in_7_14_port, 
      sum_B_in_7_13_port, sum_B_in_7_12_port, sum_B_in_7_11_port, 
      sum_B_in_7_10_port, sum_B_in_7_9_port, sum_B_in_7_8_port, 
      sum_B_in_7_7_port, sum_B_in_7_6_port, sum_B_in_7_5_port, 
      sum_B_in_7_4_port, sum_B_in_7_3_port, sum_B_in_7_2_port, 
      sum_B_in_7_1_port, sum_B_in_7_0_port, sum_out_1_19_port, 
      sum_out_1_18_port, sum_out_1_17_port, sum_out_1_16_port, 
      sum_out_1_15_port, sum_out_1_14_port, sum_out_1_13_port, 
      sum_out_1_12_port, sum_out_1_11_port, sum_out_1_10_port, sum_out_1_9_port
      , sum_out_1_8_port, sum_out_1_7_port, sum_out_1_6_port, sum_out_1_5_port,
      sum_out_1_4_port, sum_out_1_3_port, sum_out_1_2_port, sum_out_1_1_port, 
      sum_out_1_0_port, sum_out_2_21_port, sum_out_2_20_port, sum_out_2_19_port
      , sum_out_2_18_port, sum_out_2_17_port, sum_out_2_16_port, 
      sum_out_2_15_port, sum_out_2_14_port, sum_out_2_13_port, 
      sum_out_2_12_port, sum_out_2_11_port, sum_out_2_10_port, sum_out_2_9_port
      , sum_out_2_8_port, sum_out_2_7_port, sum_out_2_6_port, sum_out_2_5_port,
      sum_out_2_4_port, sum_out_2_3_port, sum_out_2_2_port, sum_out_2_1_port, 
      sum_out_2_0_port, sum_out_3_23_port, sum_out_3_22_port, sum_out_3_21_port
      , sum_out_3_20_port, sum_out_3_19_port, sum_out_3_18_port, 
      sum_out_3_17_port, sum_out_3_16_port, sum_out_3_15_port, 
      sum_out_3_14_port, sum_out_3_13_port, sum_out_3_12_port, 
      sum_out_3_11_port, sum_out_3_10_port, sum_out_3_9_port, sum_out_3_8_port,
      sum_out_3_7_port, sum_out_3_6_port, sum_out_3_5_port, sum_out_3_4_port, 
      sum_out_3_3_port, sum_out_3_2_port, sum_out_3_1_port, sum_out_3_0_port, 
      sum_out_4_25_port, sum_out_4_24_port, sum_out_4_23_port, 
      sum_out_4_22_port, sum_out_4_21_port, sum_out_4_20_port, 
      sum_out_4_19_port, sum_out_4_18_port, sum_out_4_17_port, 
      sum_out_4_16_port, sum_out_4_15_port, sum_out_4_14_port, 
      sum_out_4_13_port, sum_out_4_12_port, sum_out_4_11_port, 
      sum_out_4_10_port, sum_out_4_9_port, sum_out_4_8_port, sum_out_4_7_port, 
      sum_out_4_6_port, sum_out_4_5_port, sum_out_4_4_port, sum_out_4_3_port, 
      sum_out_4_2_port, sum_out_4_1_port, sum_out_4_0_port, sum_out_5_27_port, 
      sum_out_5_26_port, sum_out_5_25_port, sum_out_5_24_port, 
      sum_out_5_23_port, sum_out_5_22_port, sum_out_5_21_port, 
      sum_out_5_20_port, sum_out_5_19_port, sum_out_5_18_port, 
      sum_out_5_17_port, sum_out_5_16_port, sum_out_5_15_port, 
      sum_out_5_14_port, sum_out_5_13_port, sum_out_5_12_port, 
      sum_out_5_11_port, sum_out_5_10_port, sum_out_5_9_port, sum_out_5_8_port,
      sum_out_5_7_port, sum_out_5_6_port, sum_out_5_5_port, sum_out_5_4_port, 
      sum_out_5_3_port, sum_out_5_2_port, sum_out_5_1_port, sum_out_5_0_port, 
      sum_out_6_29_port, sum_out_6_28_port, sum_out_6_27_port, 
      sum_out_6_26_port, sum_out_6_25_port, sum_out_6_24_port, 
      sum_out_6_23_port, sum_out_6_22_port, sum_out_6_21_port, 
      sum_out_6_20_port, sum_out_6_19_port, sum_out_6_18_port, 
      sum_out_6_17_port, sum_out_6_16_port, sum_out_6_15_port, 
      sum_out_6_14_port, sum_out_6_13_port, sum_out_6_12_port, 
      sum_out_6_11_port, sum_out_6_10_port, sum_out_6_9_port, sum_out_6_8_port,
      sum_out_6_7_port, sum_out_6_6_port, sum_out_6_5_port, sum_out_6_4_port, 
      sum_out_6_3_port, sum_out_6_2_port, sum_out_6_1_port, sum_out_6_0_port, 
      muxes_in_3_23_port, muxes_in_3_24_port, muxes_in_3_25_port, 
      muxes_in_3_26_port, muxes_in_3_27_port, muxes_in_3_28_port, 
      muxes_in_3_29_port, muxes_in_3_30_port, muxes_in_3_31_port, 
      muxes_in_3_32_port, muxes_in_3_33_port, muxes_in_3_34_port, 
      muxes_in_3_35_port, muxes_in_3_36_port, muxes_in_3_37_port, 
      muxes_in_3_38_port, muxes_in_3_39_port, muxes_in_3_40_port, 
      muxes_in_3_41_port, muxes_in_3_42_port, muxes_in_3_43_port, 
      muxes_in_3_46_port, muxes_in_3_47_port, muxes_in_3_48_port, 
      muxes_in_3_49_port, muxes_in_3_50_port, muxes_in_3_51_port, 
      muxes_in_3_52_port, muxes_in_3_53_port, muxes_in_3_54_port, 
      muxes_in_3_55_port, muxes_in_3_56_port, muxes_in_3_57_port, 
      muxes_in_3_58_port, muxes_in_3_59_port, muxes_in_3_60_port, 
      muxes_in_3_61_port, muxes_in_3_62_port, muxes_in_3_63_port, 
      muxes_in_3_64_port, muxes_in_3_65_port, muxes_in_3_66_port, 
      muxes_in_3_138_port, muxes_in_3_139_port, muxes_in_3_140_port, 
      muxes_in_3_141_port, muxes_in_3_142_port, muxes_in_3_143_port, 
      muxes_in_3_144_port, muxes_in_3_145_port, muxes_in_3_146_port, 
      muxes_in_3_147_port, muxes_in_3_148_port, muxes_in_3_149_port, 
      muxes_in_3_150_port, muxes_in_3_151_port, muxes_in_3_152_port, 
      muxes_in_3_153_port, muxes_in_3_154_port, muxes_in_3_155_port, 
      muxes_in_3_156_port, muxes_in_3_157_port, muxes_in_3_158_port, 
      muxes_in_3_161_port, muxes_in_3_162_port, muxes_in_3_163_port, 
      muxes_in_3_164_port, muxes_in_3_165_port, muxes_in_3_166_port, 
      muxes_in_3_167_port, muxes_in_3_168_port, muxes_in_3_169_port, 
      muxes_in_3_170_port, muxes_in_3_171_port, muxes_in_3_172_port, 
      muxes_in_3_173_port, muxes_in_3_174_port, muxes_in_3_175_port, 
      muxes_in_3_176_port, muxes_in_3_177_port, muxes_in_3_178_port, 
      muxes_in_3_179_port, muxes_in_3_180_port, muxes_in_3_181_port, 
      muxes_in_4_25_port, muxes_in_4_26_port, muxes_in_4_27_port, 
      muxes_in_4_28_port, muxes_in_4_29_port, muxes_in_4_30_port, 
      muxes_in_4_31_port, muxes_in_4_32_port, muxes_in_4_33_port, 
      muxes_in_4_34_port, muxes_in_4_35_port, muxes_in_4_36_port, 
      muxes_in_4_37_port, muxes_in_4_38_port, muxes_in_4_39_port, 
      muxes_in_4_40_port, muxes_in_4_41_port, muxes_in_4_42_port, 
      muxes_in_4_43_port, muxes_in_4_44_port, muxes_in_4_45_port, 
      muxes_in_4_46_port, muxes_in_4_47_port, muxes_in_4_50_port, 
      muxes_in_4_51_port, muxes_in_4_52_port, muxes_in_4_53_port, 
      muxes_in_4_54_port, muxes_in_4_55_port, muxes_in_4_56_port, 
      muxes_in_4_57_port, muxes_in_4_58_port, muxes_in_4_59_port, 
      muxes_in_4_60_port, muxes_in_4_61_port, muxes_in_4_62_port, 
      muxes_in_4_63_port, muxes_in_4_64_port, muxes_in_4_65_port, 
      muxes_in_4_66_port, muxes_in_4_67_port, muxes_in_4_68_port, 
      muxes_in_4_69_port, muxes_in_4_70_port, muxes_in_4_71_port, 
      muxes_in_4_72_port, muxes_in_4_150_port, muxes_in_4_151_port, 
      muxes_in_4_152_port, muxes_in_4_153_port, muxes_in_4_154_port, 
      muxes_in_4_155_port, muxes_in_4_156_port, muxes_in_4_157_port, 
      muxes_in_4_158_port, muxes_in_4_159_port, muxes_in_4_160_port, 
      muxes_in_4_161_port, muxes_in_4_162_port, muxes_in_4_163_port, 
      muxes_in_4_164_port, muxes_in_4_165_port, muxes_in_4_166_port, 
      muxes_in_4_167_port, muxes_in_4_168_port, muxes_in_4_169_port, 
      muxes_in_4_170_port, muxes_in_4_171_port, muxes_in_4_172_port, 
      muxes_in_4_175_port, muxes_in_4_176_port, muxes_in_4_177_port, 
      muxes_in_4_178_port, muxes_in_4_179_port, muxes_in_4_180_port, 
      muxes_in_4_181_port, muxes_in_4_182_port, muxes_in_4_183_port, 
      muxes_in_4_184_port, muxes_in_4_185_port, muxes_in_4_186_port, 
      muxes_in_4_187_port, muxes_in_4_188_port, muxes_in_4_189_port, 
      muxes_in_4_190_port, muxes_in_4_191_port, muxes_in_4_192_port, 
      muxes_in_4_193_port, muxes_in_4_194_port, muxes_in_4_195_port, 
      muxes_in_4_196_port, muxes_in_4_197_port, muxes_in_5_27_port, 
      muxes_in_5_28_port, muxes_in_5_29_port, muxes_in_5_30_port, 
      muxes_in_5_31_port, muxes_in_5_32_port, muxes_in_5_33_port, 
      muxes_in_5_34_port, muxes_in_5_35_port, muxes_in_5_36_port, 
      muxes_in_5_37_port, muxes_in_5_38_port, muxes_in_5_39_port, 
      muxes_in_5_40_port, muxes_in_5_41_port, muxes_in_5_42_port, 
      muxes_in_5_43_port, muxes_in_5_44_port, muxes_in_5_45_port, 
      muxes_in_5_46_port, muxes_in_5_47_port, muxes_in_5_48_port, 
      muxes_in_5_49_port, muxes_in_5_50_port, muxes_in_5_51_port, 
      muxes_in_5_54_port, muxes_in_5_55_port, muxes_in_5_56_port, 
      muxes_in_5_57_port, muxes_in_5_58_port, muxes_in_5_59_port, 
      muxes_in_5_60_port, muxes_in_5_61_port, muxes_in_5_62_port, 
      muxes_in_5_63_port, muxes_in_5_64_port, muxes_in_5_65_port, 
      muxes_in_5_66_port, muxes_in_5_67_port, muxes_in_5_68_port, 
      muxes_in_5_69_port, muxes_in_5_70_port, muxes_in_5_71_port, 
      muxes_in_5_72_port, muxes_in_5_73_port, muxes_in_5_74_port, 
      muxes_in_5_75_port, muxes_in_5_76_port, muxes_in_5_77_port, 
      muxes_in_5_78_port, muxes_in_5_162_port, muxes_in_5_163_port, 
      muxes_in_5_164_port, muxes_in_5_165_port, muxes_in_5_166_port, 
      muxes_in_5_167_port, muxes_in_5_168_port, muxes_in_5_169_port, 
      muxes_in_5_170_port, muxes_in_5_171_port, muxes_in_5_172_port, 
      muxes_in_5_173_port, muxes_in_5_174_port, muxes_in_5_175_port, 
      muxes_in_5_176_port, muxes_in_5_177_port, muxes_in_5_178_port, 
      muxes_in_5_179_port, muxes_in_5_180_port, muxes_in_5_181_port, 
      muxes_in_5_182_port, muxes_in_5_183_port, muxes_in_5_184_port, 
      muxes_in_5_185_port, muxes_in_5_186_port, muxes_in_5_189_port, 
      muxes_in_5_190_port, muxes_in_5_191_port, muxes_in_5_192_port, 
      muxes_in_5_193_port, muxes_in_5_194_port, muxes_in_5_195_port, 
      muxes_in_5_196_port, muxes_in_5_197_port, muxes_in_5_198_port, 
      muxes_in_5_199_port, muxes_in_5_200_port, muxes_in_5_201_port, 
      muxes_in_5_202_port, muxes_in_5_203_port, muxes_in_5_204_port, 
      muxes_in_5_205_port, muxes_in_5_206_port, muxes_in_5_207_port, 
      muxes_in_5_208_port, muxes_in_5_209_port, muxes_in_5_210_port, 
      muxes_in_5_211_port, muxes_in_5_212_port, muxes_in_5_213_port, 
      muxes_in_6_29_port, muxes_in_6_30_port, muxes_in_6_31_port, 
      muxes_in_6_32_port, muxes_in_6_33_port, muxes_in_6_34_port, 
      muxes_in_6_35_port, muxes_in_6_36_port, muxes_in_6_37_port, 
      muxes_in_6_38_port, muxes_in_6_39_port, muxes_in_6_40_port, 
      muxes_in_6_41_port, muxes_in_6_42_port, muxes_in_6_43_port, 
      muxes_in_6_44_port, muxes_in_6_45_port, muxes_in_6_46_port, 
      muxes_in_6_47_port, muxes_in_6_48_port, muxes_in_6_49_port, 
      muxes_in_6_50_port, muxes_in_6_51_port, muxes_in_6_52_port, 
      muxes_in_6_53_port, muxes_in_6_54_port, muxes_in_6_55_port, 
      muxes_in_6_58_port, muxes_in_6_59_port, muxes_in_6_60_port, 
      muxes_in_6_61_port, muxes_in_6_62_port, muxes_in_6_63_port, 
      muxes_in_6_64_port, muxes_in_6_65_port, muxes_in_6_66_port, 
      muxes_in_6_67_port, muxes_in_6_68_port, muxes_in_6_69_port, 
      muxes_in_6_70_port, muxes_in_6_71_port, muxes_in_6_72_port, 
      muxes_in_6_73_port, muxes_in_6_74_port, muxes_in_6_75_port, 
      muxes_in_6_76_port, muxes_in_6_77_port, muxes_in_6_78_port, 
      muxes_in_6_79_port, muxes_in_6_80_port, muxes_in_6_81_port, 
      muxes_in_6_82_port, muxes_in_6_83_port, muxes_in_6_84_port, 
      muxes_in_6_174_port, muxes_in_6_175_port, muxes_in_6_176_port, 
      muxes_in_6_177_port, muxes_in_6_178_port, muxes_in_6_179_port, 
      muxes_in_6_180_port, muxes_in_6_181_port, muxes_in_6_182_port, 
      muxes_in_6_183_port, muxes_in_6_184_port, muxes_in_6_185_port, 
      muxes_in_6_186_port, muxes_in_6_187_port, muxes_in_6_188_port, 
      muxes_in_6_189_port, muxes_in_6_190_port, muxes_in_6_191_port, 
      muxes_in_6_192_port, muxes_in_6_193_port, muxes_in_6_194_port, 
      muxes_in_6_195_port, muxes_in_6_196_port, muxes_in_6_197_port, 
      muxes_in_6_198_port, muxes_in_6_199_port, muxes_in_6_200_port, 
      muxes_in_6_203_port, muxes_in_6_204_port, muxes_in_6_205_port, 
      muxes_in_6_206_port, muxes_in_6_207_port, muxes_in_6_208_port, 
      muxes_in_6_209_port, muxes_in_6_210_port, muxes_in_6_211_port, 
      muxes_in_6_212_port, muxes_in_6_213_port, muxes_in_6_214_port, 
      muxes_in_6_215_port, muxes_in_6_216_port, muxes_in_6_217_port, 
      muxes_in_6_218_port, muxes_in_6_219_port, muxes_in_6_220_port, 
      muxes_in_6_221_port, muxes_in_6_222_port, muxes_in_6_223_port, 
      muxes_in_6_224_port, muxes_in_6_225_port, muxes_in_6_226_port, 
      muxes_in_6_227_port, muxes_in_6_228_port, muxes_in_6_229_port, 
      muxes_in_7_31_port, muxes_in_7_32_port, muxes_in_7_33_port, 
      muxes_in_7_34_port, muxes_in_7_35_port, muxes_in_7_36_port, 
      muxes_in_7_37_port, muxes_in_7_38_port, muxes_in_7_39_port, 
      muxes_in_7_40_port, muxes_in_7_41_port, muxes_in_7_42_port, 
      muxes_in_7_43_port, muxes_in_7_44_port, muxes_in_7_45_port, 
      muxes_in_7_46_port, muxes_in_7_47_port, muxes_in_7_48_port, 
      muxes_in_7_49_port, muxes_in_7_50_port, muxes_in_7_51_port, 
      muxes_in_7_52_port, muxes_in_7_53_port, muxes_in_7_54_port, 
      muxes_in_7_55_port, muxes_in_7_56_port, muxes_in_7_57_port, 
      muxes_in_7_58_port, muxes_in_7_59_port, muxes_in_7_62_port, 
      muxes_in_7_63_port, muxes_in_7_64_port, muxes_in_7_65_port, 
      muxes_in_7_66_port, muxes_in_7_67_port, muxes_in_7_68_port, 
      muxes_in_7_69_port, muxes_in_7_70_port, muxes_in_7_71_port, 
      muxes_in_7_72_port, muxes_in_7_73_port, muxes_in_7_74_port, 
      muxes_in_7_75_port, muxes_in_7_76_port, muxes_in_7_77_port, 
      muxes_in_7_78_port, muxes_in_7_79_port, muxes_in_7_80_port, 
      muxes_in_7_81_port, muxes_in_7_82_port, muxes_in_7_83_port, 
      muxes_in_7_84_port, muxes_in_7_85_port, muxes_in_7_86_port, 
      muxes_in_7_87_port, muxes_in_7_88_port, muxes_in_7_89_port, 
      muxes_in_7_90_port, muxes_in_7_186_port, muxes_in_7_187_port, 
      muxes_in_7_188_port, muxes_in_7_189_port, muxes_in_7_190_port, 
      muxes_in_7_191_port, muxes_in_7_192_port, muxes_in_7_193_port, 
      muxes_in_7_194_port, muxes_in_7_195_port, muxes_in_7_196_port, 
      muxes_in_7_197_port, muxes_in_7_198_port, muxes_in_7_199_port, 
      muxes_in_7_200_port, muxes_in_7_201_port, muxes_in_7_202_port, 
      muxes_in_7_203_port, muxes_in_7_204_port, muxes_in_7_205_port, 
      muxes_in_7_206_port, muxes_in_7_207_port, muxes_in_7_208_port, 
      muxes_in_7_209_port, muxes_in_7_210_port, muxes_in_7_211_port, 
      muxes_in_7_212_port, muxes_in_7_213_port, muxes_in_7_214_port, 
      muxes_in_7_217_port, muxes_in_7_218_port, muxes_in_7_219_port, 
      muxes_in_7_220_port, muxes_in_7_221_port, muxes_in_7_222_port, 
      muxes_in_7_223_port, muxes_in_7_224_port, muxes_in_7_225_port, 
      muxes_in_7_226_port, muxes_in_7_227_port, muxes_in_7_228_port, 
      muxes_in_7_229_port, muxes_in_7_230_port, muxes_in_7_231_port, 
      muxes_in_7_232_port, muxes_in_7_233_port, muxes_in_7_234_port, 
      muxes_in_7_235_port, muxes_in_7_236_port, muxes_in_7_237_port, 
      muxes_in_7_238_port, muxes_in_7_239_port, muxes_in_7_240_port, 
      muxes_in_7_241_port, muxes_in_7_242_port, muxes_in_7_243_port, 
      muxes_in_7_244_port, muxes_in_7_245_port, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363
      , n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372,
      n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, 
      n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, 
      n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, 
      n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, 
      n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, 
      n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, 
      n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, 
      n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, 
      n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, 
      n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, 
      n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, 
      n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, 
      n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, 
      n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, 
      n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, 
      n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, 
      n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, 
      n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, 
      n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, 
      n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, 
      n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, 
      n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, 
      n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, 
      n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, 
      n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, 
      n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, 
      n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, 
      n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, 
      n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, 
      n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, 
      n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, 
      n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, 
      n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, 
      n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, 
      n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, 
      n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, 
      n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, 
      n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, 
      n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, 
      n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, 
      n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, 
      n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, 
      n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, 
      n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, 
      n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, 
      n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, 
      n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, 
      n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, 
      n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, 
      n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, 
      n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, 
      n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, 
      n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, 
      n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, 
      n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, 
      n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, 
      n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, 
      n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, 
      n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, 
      n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, 
      n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, 
      n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, 
      n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, 
      n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, 
      n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, 
      n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, 
      n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, 
      n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, 
      n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, 
      n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, 
      n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, 
      n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, 
      n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, 
      n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, 
      n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, 
      n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, 
      n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, 
      n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, 
      n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, 
      n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, 
      n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, 
      n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, 
      n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, 
      n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, 
      n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, 
      n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, 
      n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, 
      n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, 
      n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, 
      n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, 
      n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, 
      n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, 
      n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, 
      n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, 
      n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, 
      n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, 
      n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, 
      n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, 
      n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, 
      n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, 
      n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, 
      n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, 
      n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, 
      n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, 
      n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, 
      n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, 
      n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, 
      n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, 
      n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, 
      n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, 
      n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, 
      n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, 
      n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, 
      n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, 
      n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, 
      n_4408, n_4409, n_4410, n_4411 : std_logic;

begin
   
   X_Logic0_port <= '0';
   minusA_0 : complement2_N17 port map( value_in(16) => multiplier(15), 
                           value_in(15) => multiplier(15), value_in(14) => 
                           multiplier(14), value_in(13) => multiplier(13), 
                           value_in(12) => multiplier(12), value_in(11) => 
                           multiplier(11), value_in(10) => multiplier(10), 
                           value_in(9) => multiplier(9), value_in(8) => 
                           multiplier(8), value_in(7) => multiplier(7), 
                           value_in(6) => multiplier(6), value_in(5) => 
                           multiplier(5), value_in(4) => multiplier(4), 
                           value_in(3) => multiplier(3), value_in(2) => 
                           multiplier(2), value_in(1) => multiplier(1), 
                           value_in(0) => multiplier(0), value_out(16) => 
                           muxes_in_0_119_port, value_out(15) => 
                           muxes_in_0_102_port, value_out(14) => 
                           muxes_in_0_103_port, value_out(13) => 
                           muxes_in_0_104_port, value_out(12) => 
                           muxes_in_0_105_port, value_out(11) => 
                           muxes_in_0_106_port, value_out(10) => 
                           muxes_in_0_107_port, value_out(9) => 
                           muxes_in_0_108_port, value_out(8) => 
                           muxes_in_0_109_port, value_out(7) => 
                           muxes_in_0_110_port, value_out(6) => 
                           muxes_in_0_111_port, value_out(5) => 
                           muxes_in_0_112_port, value_out(4) => 
                           muxes_in_0_113_port, value_out(3) => 
                           muxes_in_0_114_port, value_out(2) => 
                           muxes_in_0_115_port, value_out(1) => 
                           muxes_in_0_116_port, value_out(0) => 
                           muxes_in_0_117_port);
   ENC0_0 : encoder_0 port map( y(2) => multiplicand(1), y(1) => 
                           multiplicand(0), y(0) => X_Logic0_port, sel(2) => 
                           encoder_out_0_2_port, sel(1) => encoder_out_0_1_port
                           , sel(0) => encoder_out_0_0_port);
   MUX0_0 : MUX_zbit_nbit_N17_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => multiplier(15), inputs(18) => 
                           multiplier(15), inputs(19) => multiplier(14), 
                           inputs(20) => multiplier(13), inputs(21) => 
                           multiplier(12), inputs(22) => multiplier(11), 
                           inputs(23) => multiplier(10), inputs(24) => 
                           multiplier(9), inputs(25) => multiplier(8), 
                           inputs(26) => multiplier(7), inputs(27) => 
                           multiplier(6), inputs(28) => multiplier(5), 
                           inputs(29) => multiplier(4), inputs(30) => 
                           multiplier(3), inputs(31) => multiplier(2), 
                           inputs(32) => multiplier(1), inputs(33) => 
                           multiplier(0), inputs(34) => multiplier(15), 
                           inputs(35) => multiplier(14), inputs(36) => 
                           multiplier(13), inputs(37) => multiplier(12), 
                           inputs(38) => multiplier(11), inputs(39) => 
                           multiplier(10), inputs(40) => multiplier(9), 
                           inputs(41) => multiplier(8), inputs(42) => 
                           multiplier(7), inputs(43) => multiplier(6), 
                           inputs(44) => multiplier(5), inputs(45) => 
                           multiplier(4), inputs(46) => multiplier(3), 
                           inputs(47) => multiplier(2), inputs(48) => 
                           multiplier(1), inputs(49) => multiplier(0), 
                           inputs(50) => X_Logic0_port, inputs(51) => 
                           X_Logic0_port, inputs(52) => X_Logic0_port, 
                           inputs(53) => X_Logic0_port, inputs(54) => 
                           X_Logic0_port, inputs(55) => X_Logic0_port, 
                           inputs(56) => X_Logic0_port, inputs(57) => 
                           X_Logic0_port, inputs(58) => X_Logic0_port, 
                           inputs(59) => X_Logic0_port, inputs(60) => 
                           X_Logic0_port, inputs(61) => X_Logic0_port, 
                           inputs(62) => X_Logic0_port, inputs(63) => 
                           X_Logic0_port, inputs(64) => X_Logic0_port, 
                           inputs(65) => X_Logic0_port, inputs(66) => 
                           X_Logic0_port, inputs(67) => X_Logic0_port, 
                           inputs(68) => X_Logic0_port, inputs(69) => 
                           X_Logic0_port, inputs(70) => X_Logic0_port, 
                           inputs(71) => X_Logic0_port, inputs(72) => 
                           X_Logic0_port, inputs(73) => X_Logic0_port, 
                           inputs(74) => X_Logic0_port, inputs(75) => 
                           X_Logic0_port, inputs(76) => X_Logic0_port, 
                           inputs(77) => X_Logic0_port, inputs(78) => 
                           X_Logic0_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           muxes_in_0_102_port, inputs(103) => 
                           muxes_in_0_103_port, inputs(104) => 
                           muxes_in_0_104_port, inputs(105) => 
                           muxes_in_0_105_port, inputs(106) => 
                           muxes_in_0_106_port, inputs(107) => 
                           muxes_in_0_107_port, inputs(108) => 
                           muxes_in_0_108_port, inputs(109) => 
                           muxes_in_0_109_port, inputs(110) => 
                           muxes_in_0_110_port, inputs(111) => 
                           muxes_in_0_111_port, inputs(112) => 
                           muxes_in_0_112_port, inputs(113) => 
                           muxes_in_0_113_port, inputs(114) => 
                           muxes_in_0_114_port, inputs(115) => 
                           muxes_in_0_115_port, inputs(116) => 
                           muxes_in_0_116_port, inputs(117) => 
                           muxes_in_0_117_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => muxes_in_0_119_port, inputs(120) => 
                           muxes_in_0_102_port, inputs(121) => 
                           muxes_in_0_103_port, inputs(122) => 
                           muxes_in_0_104_port, inputs(123) => 
                           muxes_in_0_105_port, inputs(124) => 
                           muxes_in_0_106_port, inputs(125) => 
                           muxes_in_0_107_port, inputs(126) => 
                           muxes_in_0_108_port, inputs(127) => 
                           muxes_in_0_109_port, inputs(128) => 
                           muxes_in_0_110_port, inputs(129) => 
                           muxes_in_0_111_port, inputs(130) => 
                           muxes_in_0_112_port, inputs(131) => 
                           muxes_in_0_113_port, inputs(132) => 
                           muxes_in_0_114_port, inputs(133) => 
                           muxes_in_0_115_port, inputs(134) => 
                           muxes_in_0_116_port, inputs(135) => 
                           muxes_in_0_117_port, SEL(2) => encoder_out_0_2_port,
                           SEL(1) => encoder_out_0_1_port, SEL(0) => 
                           encoder_out_0_0_port, Y(16) => sum_B_in_1_18_port, 
                           Y(15) => sum_B_in_1_15_port, Y(14) => 
                           sum_B_in_1_14_port, Y(13) => sum_B_in_1_13_port, 
                           Y(12) => sum_B_in_1_12_port, Y(11) => 
                           sum_B_in_1_11_port, Y(10) => sum_B_in_1_10_port, 
                           Y(9) => sum_B_in_1_9_port, Y(8) => sum_B_in_1_8_port
                           , Y(7) => sum_B_in_1_7_port, Y(6) => 
                           sum_B_in_1_6_port, Y(5) => sum_B_in_1_5_port, Y(4) 
                           => sum_B_in_1_4_port, Y(3) => sum_B_in_1_3_port, 
                           Y(2) => sum_B_in_1_2_port, Y(1) => sum_B_in_1_1_port
                           , Y(0) => sum_B_in_1_0_port);
   ENCi_1 : encoder_7 port map( y(2) => multiplicand(3), y(1) => 
                           multiplicand(2), y(0) => multiplicand(1), sel(2) => 
                           encoder_out_1_2_port, sel(1) => encoder_out_1_1_port
                           , sel(0) => encoder_out_1_0_port);
   MUXi_1 : MUX_zbit_nbit_N19_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => multiplier(15), 
                           inputs(20) => multiplier(15), inputs(21) => 
                           multiplier(14), inputs(22) => multiplier(13), 
                           inputs(23) => multiplier(12), inputs(24) => 
                           multiplier(11), inputs(25) => multiplier(10), 
                           inputs(26) => multiplier(9), inputs(27) => 
                           multiplier(8), inputs(28) => multiplier(7), 
                           inputs(29) => multiplier(6), inputs(30) => 
                           multiplier(5), inputs(31) => multiplier(4), 
                           inputs(32) => multiplier(3), inputs(33) => 
                           multiplier(2), inputs(34) => multiplier(1), 
                           inputs(35) => multiplier(0), inputs(36) => 
                           X_Logic0_port, inputs(37) => X_Logic0_port, 
                           inputs(38) => multiplier(15), inputs(39) => 
                           multiplier(14), inputs(40) => multiplier(13), 
                           inputs(41) => multiplier(12), inputs(42) => 
                           multiplier(11), inputs(43) => multiplier(10), 
                           inputs(44) => multiplier(9), inputs(45) => 
                           multiplier(8), inputs(46) => multiplier(7), 
                           inputs(47) => multiplier(6), inputs(48) => 
                           multiplier(5), inputs(49) => multiplier(4), 
                           inputs(50) => multiplier(3), inputs(51) => 
                           multiplier(2), inputs(52) => multiplier(1), 
                           inputs(53) => multiplier(0), inputs(54) => 
                           X_Logic0_port, inputs(55) => X_Logic0_port, 
                           inputs(56) => X_Logic0_port, inputs(57) => 
                           X_Logic0_port, inputs(58) => X_Logic0_port, 
                           inputs(59) => X_Logic0_port, inputs(60) => 
                           X_Logic0_port, inputs(61) => X_Logic0_port, 
                           inputs(62) => X_Logic0_port, inputs(63) => 
                           X_Logic0_port, inputs(64) => X_Logic0_port, 
                           inputs(65) => X_Logic0_port, inputs(66) => 
                           X_Logic0_port, inputs(67) => X_Logic0_port, 
                           inputs(68) => X_Logic0_port, inputs(69) => 
                           X_Logic0_port, inputs(70) => X_Logic0_port, 
                           inputs(71) => X_Logic0_port, inputs(72) => 
                           X_Logic0_port, inputs(73) => X_Logic0_port, 
                           inputs(74) => X_Logic0_port, inputs(75) => 
                           X_Logic0_port, inputs(76) => X_Logic0_port, 
                           inputs(77) => X_Logic0_port, inputs(78) => 
                           X_Logic0_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           muxes_in_0_102_port, inputs(115) => 
                           muxes_in_0_103_port, inputs(116) => 
                           muxes_in_0_104_port, inputs(117) => 
                           muxes_in_0_105_port, inputs(118) => 
                           muxes_in_0_106_port, inputs(119) => 
                           muxes_in_0_107_port, inputs(120) => 
                           muxes_in_0_108_port, inputs(121) => 
                           muxes_in_0_109_port, inputs(122) => 
                           muxes_in_0_110_port, inputs(123) => 
                           muxes_in_0_111_port, inputs(124) => 
                           muxes_in_0_112_port, inputs(125) => 
                           muxes_in_0_113_port, inputs(126) => 
                           muxes_in_0_114_port, inputs(127) => 
                           muxes_in_0_115_port, inputs(128) => 
                           muxes_in_0_116_port, inputs(129) => 
                           muxes_in_0_117_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => muxes_in_0_119_port, 
                           inputs(134) => muxes_in_0_102_port, inputs(135) => 
                           muxes_in_0_103_port, inputs(136) => 
                           muxes_in_0_104_port, inputs(137) => 
                           muxes_in_0_105_port, inputs(138) => 
                           muxes_in_0_106_port, inputs(139) => 
                           muxes_in_0_107_port, inputs(140) => 
                           muxes_in_0_108_port, inputs(141) => 
                           muxes_in_0_109_port, inputs(142) => 
                           muxes_in_0_110_port, inputs(143) => 
                           muxes_in_0_111_port, inputs(144) => 
                           muxes_in_0_112_port, inputs(145) => 
                           muxes_in_0_113_port, inputs(146) => 
                           muxes_in_0_114_port, inputs(147) => 
                           muxes_in_0_115_port, inputs(148) => 
                           muxes_in_0_116_port, inputs(149) => 
                           muxes_in_0_117_port, inputs(150) => X_Logic0_port, 
                           inputs(151) => X_Logic0_port, SEL(2) => 
                           encoder_out_1_2_port, SEL(1) => encoder_out_1_1_port
                           , SEL(0) => encoder_out_1_0_port, Y(18) => 
                           mux_out_1_18_port, Y(17) => mux_out_1_17_port, Y(16)
                           => mux_out_1_16_port, Y(15) => mux_out_1_15_port, 
                           Y(14) => mux_out_1_14_port, Y(13) => 
                           mux_out_1_13_port, Y(12) => mux_out_1_12_port, Y(11)
                           => mux_out_1_11_port, Y(10) => mux_out_1_10_port, 
                           Y(9) => mux_out_1_9_port, Y(8) => mux_out_1_8_port, 
                           Y(7) => mux_out_1_7_port, Y(6) => mux_out_1_6_port, 
                           Y(5) => mux_out_1_5_port, Y(4) => mux_out_1_4_port, 
                           Y(3) => mux_out_1_3_port, Y(2) => mux_out_1_2_port, 
                           Y(1) => mux_out_1_1_port, Y(0) => mux_out_1_0_port);
   ADD1_1 : adder_NBIT19 port map( a(18) => mux_out_1_18_port, a(17) => 
                           mux_out_1_17_port, a(16) => mux_out_1_16_port, a(15)
                           => mux_out_1_15_port, a(14) => mux_out_1_14_port, 
                           a(13) => mux_out_1_13_port, a(12) => 
                           mux_out_1_12_port, a(11) => mux_out_1_11_port, a(10)
                           => mux_out_1_10_port, a(9) => mux_out_1_9_port, a(8)
                           => mux_out_1_8_port, a(7) => mux_out_1_7_port, a(6) 
                           => mux_out_1_6_port, a(5) => mux_out_1_5_port, a(4) 
                           => mux_out_1_4_port, a(3) => mux_out_1_3_port, a(2) 
                           => mux_out_1_2_port, a(1) => mux_out_1_1_port, a(0) 
                           => mux_out_1_0_port, b(18) => sum_B_in_1_18_port, 
                           b(17) => sum_B_in_1_18_port, b(16) => 
                           sum_B_in_1_18_port, b(15) => sum_B_in_1_15_port, 
                           b(14) => sum_B_in_1_14_port, b(13) => 
                           sum_B_in_1_13_port, b(12) => sum_B_in_1_12_port, 
                           b(11) => sum_B_in_1_11_port, b(10) => 
                           sum_B_in_1_10_port, b(9) => sum_B_in_1_9_port, b(8) 
                           => sum_B_in_1_8_port, b(7) => sum_B_in_1_7_port, 
                           b(6) => sum_B_in_1_6_port, b(5) => sum_B_in_1_5_port
                           , b(4) => sum_B_in_1_4_port, b(3) => 
                           sum_B_in_1_3_port, b(2) => sum_B_in_1_2_port, b(1) 
                           => sum_B_in_1_1_port, b(0) => sum_B_in_1_0_port, cin
                           => X_Logic0_port, s(19) => sum_out_1_19_port, s(18) 
                           => sum_out_1_18_port, s(17) => sum_out_1_17_port, 
                           s(16) => sum_out_1_16_port, s(15) => 
                           sum_out_1_15_port, s(14) => sum_out_1_14_port, s(13)
                           => sum_out_1_13_port, s(12) => sum_out_1_12_port, 
                           s(11) => sum_out_1_11_port, s(10) => 
                           sum_out_1_10_port, s(9) => sum_out_1_9_port, s(8) =>
                           sum_out_1_8_port, s(7) => sum_out_1_7_port, s(6) => 
                           sum_out_1_6_port, s(5) => sum_out_1_5_port, s(4) => 
                           sum_out_1_4_port, s(3) => sum_out_1_3_port, s(2) => 
                           sum_out_1_2_port, s(1) => sum_out_1_1_port, s(0) => 
                           sum_out_1_0_port);
   pip_del_reg_add1_1 : reg_nbit_n32_6 port map( clk => n12, reset => n5, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           X_Logic0_port, d(20) => X_Logic0_port, d(19) => 
                           sum_out_1_19_port, d(18) => sum_out_1_18_port, d(17)
                           => sum_out_1_17_port, d(16) => sum_out_1_16_port, 
                           d(15) => sum_out_1_15_port, d(14) => 
                           sum_out_1_14_port, d(13) => sum_out_1_13_port, d(12)
                           => sum_out_1_12_port, d(11) => sum_out_1_11_port, 
                           d(10) => sum_out_1_10_port, d(9) => sum_out_1_9_port
                           , d(8) => sum_out_1_8_port, d(7) => sum_out_1_7_port
                           , d(6) => sum_out_1_6_port, d(5) => sum_out_1_5_port
                           , d(4) => sum_out_1_4_port, d(3) => sum_out_1_3_port
                           , d(2) => sum_out_1_2_port, d(1) => sum_out_1_1_port
                           , d(0) => sum_out_1_0_port, Q(31) => n_3357, Q(30) 
                           => n_3358, Q(29) => n_3359, Q(28) => n_3360, Q(27) 
                           => n_3361, Q(26) => n_3362, Q(25) => n_3363, Q(24) 
                           => n_3364, Q(23) => n_3365, Q(22) => n_3366, Q(21) 
                           => n_3367, Q(20) => n_3368, Q(19) => n_3369, Q(18) 
                           => sum_B_in_2_20_port, Q(17) => sum_B_in_2_17_port, 
                           Q(16) => sum_B_in_2_16_port, Q(15) => 
                           sum_B_in_2_15_port, Q(14) => sum_B_in_2_14_port, 
                           Q(13) => sum_B_in_2_13_port, Q(12) => 
                           sum_B_in_2_12_port, Q(11) => sum_B_in_2_11_port, 
                           Q(10) => sum_B_in_2_10_port, Q(9) => 
                           sum_B_in_2_9_port, Q(8) => sum_B_in_2_8_port, Q(7) 
                           => sum_B_in_2_7_port, Q(6) => sum_B_in_2_6_port, 
                           Q(5) => sum_B_in_2_5_port, Q(4) => sum_B_in_2_4_port
                           , Q(3) => sum_B_in_2_3_port, Q(2) => 
                           sum_B_in_2_2_port, Q(1) => sum_B_in_2_1_port, Q(0) 
                           => sum_B_in_2_0_port);
   ENCi_2 : encoder_6 port map( y(2) => multiplicand_pip_2_5_port, y(1) => 
                           multiplicand_pip_2_4_port, y(0) => 
                           multiplicand_pip_2_3_port, sel(2) => 
                           encoder_out_2_2_port, sel(1) => encoder_out_2_1_port
                           , sel(0) => encoder_out_2_0_port);
   pip_del_reg_muxi_2 : reg_nbit_n249_0 port map( clk => n9, reset => n6, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => multiplier(15), 
                           d(226) => multiplier(15), d(225) => multiplier(14), 
                           d(224) => multiplier(13), d(223) => multiplier(12), 
                           d(222) => multiplier(11), d(221) => multiplier(10), 
                           d(220) => multiplier(9), d(219) => multiplier(8), 
                           d(218) => multiplier(7), d(217) => multiplier(6), 
                           d(216) => multiplier(5), d(215) => multiplier(4), 
                           d(214) => multiplier(3), d(213) => multiplier(2), 
                           d(212) => multiplier(1), d(211) => multiplier(0), 
                           d(210) => X_Logic0_port, d(209) => X_Logic0_port, 
                           d(208) => X_Logic0_port, d(207) => X_Logic0_port, 
                           d(206) => multiplier(15), d(205) => multiplier(14), 
                           d(204) => multiplier(13), d(203) => multiplier(12), 
                           d(202) => multiplier(11), d(201) => multiplier(10), 
                           d(200) => multiplier(9), d(199) => multiplier(8), 
                           d(198) => multiplier(7), d(197) => multiplier(6), 
                           d(196) => multiplier(5), d(195) => multiplier(4), 
                           d(194) => multiplier(3), d(193) => multiplier(2), 
                           d(192) => multiplier(1), d(191) => multiplier(0), 
                           d(190) => X_Logic0_port, d(189) => X_Logic0_port, 
                           d(188) => X_Logic0_port, d(187) => X_Logic0_port, 
                           d(186) => X_Logic0_port, d(185) => X_Logic0_port, 
                           d(184) => X_Logic0_port, d(183) => X_Logic0_port, 
                           d(182) => X_Logic0_port, d(181) => X_Logic0_port, 
                           d(180) => X_Logic0_port, d(179) => X_Logic0_port, 
                           d(178) => X_Logic0_port, d(177) => X_Logic0_port, 
                           d(176) => X_Logic0_port, d(175) => X_Logic0_port, 
                           d(174) => X_Logic0_port, d(173) => X_Logic0_port, 
                           d(172) => X_Logic0_port, d(171) => X_Logic0_port, 
                           d(170) => X_Logic0_port, d(169) => X_Logic0_port, 
                           d(168) => X_Logic0_port, d(167) => X_Logic0_port, 
                           d(166) => X_Logic0_port, d(165) => X_Logic0_port, 
                           d(164) => X_Logic0_port, d(163) => X_Logic0_port, 
                           d(162) => X_Logic0_port, d(161) => X_Logic0_port, 
                           d(160) => X_Logic0_port, d(159) => X_Logic0_port, 
                           d(158) => X_Logic0_port, d(157) => X_Logic0_port, 
                           d(156) => X_Logic0_port, d(155) => X_Logic0_port, 
                           d(154) => X_Logic0_port, d(153) => X_Logic0_port, 
                           d(152) => X_Logic0_port, d(151) => X_Logic0_port, 
                           d(150) => X_Logic0_port, d(149) => X_Logic0_port, 
                           d(148) => X_Logic0_port, d(147) => X_Logic0_port, 
                           d(146) => X_Logic0_port, d(145) => X_Logic0_port, 
                           d(144) => X_Logic0_port, d(143) => X_Logic0_port, 
                           d(142) => X_Logic0_port, d(141) => X_Logic0_port, 
                           d(140) => X_Logic0_port, d(139) => X_Logic0_port, 
                           d(138) => X_Logic0_port, d(137) => X_Logic0_port, 
                           d(136) => X_Logic0_port, d(135) => X_Logic0_port, 
                           d(134) => X_Logic0_port, d(133) => X_Logic0_port, 
                           d(132) => X_Logic0_port, d(131) => X_Logic0_port, 
                           d(130) => X_Logic0_port, d(129) => X_Logic0_port, 
                           d(128) => X_Logic0_port, d(127) => X_Logic0_port, 
                           d(126) => X_Logic0_port, d(125) => X_Logic0_port, 
                           d(124) => X_Logic0_port, d(123) => X_Logic0_port, 
                           d(122) => muxes_in_0_102_port, d(121) => 
                           muxes_in_0_103_port, d(120) => muxes_in_0_104_port, 
                           d(119) => muxes_in_0_105_port, d(118) => 
                           muxes_in_0_106_port, d(117) => muxes_in_0_107_port, 
                           d(116) => muxes_in_0_108_port, d(115) => 
                           muxes_in_0_109_port, d(114) => muxes_in_0_110_port, 
                           d(113) => muxes_in_0_111_port, d(112) => 
                           muxes_in_0_112_port, d(111) => muxes_in_0_113_port, 
                           d(110) => muxes_in_0_114_port, d(109) => 
                           muxes_in_0_115_port, d(108) => muxes_in_0_116_port, 
                           d(107) => muxes_in_0_117_port, d(106) => 
                           X_Logic0_port, d(105) => X_Logic0_port, d(104) => 
                           X_Logic0_port, d(103) => X_Logic0_port, d(102) => 
                           X_Logic0_port, d(101) => muxes_in_0_119_port, d(100)
                           => muxes_in_0_102_port, d(99) => muxes_in_0_103_port
                           , d(98) => muxes_in_0_104_port, d(97) => 
                           muxes_in_0_105_port, d(96) => muxes_in_0_106_port, 
                           d(95) => muxes_in_0_107_port, d(94) => 
                           muxes_in_0_108_port, d(93) => muxes_in_0_109_port, 
                           d(92) => muxes_in_0_110_port, d(91) => 
                           muxes_in_0_111_port, d(90) => muxes_in_0_112_port, 
                           d(89) => muxes_in_0_113_port, d(88) => 
                           muxes_in_0_114_port, d(87) => muxes_in_0_115_port, 
                           d(86) => muxes_in_0_116_port, d(85) => 
                           muxes_in_0_117_port, d(84) => X_Logic0_port, d(83) 
                           => X_Logic0_port, d(82) => X_Logic0_port, d(81) => 
                           X_Logic0_port, d(80) => X_Logic0_port, d(79) => 
                           X_Logic0_port, d(78) => X_Logic0_port, d(77) => 
                           X_Logic0_port, d(76) => X_Logic0_port, d(75) => 
                           X_Logic0_port, d(74) => X_Logic0_port, d(73) => 
                           X_Logic0_port, d(72) => X_Logic0_port, d(71) => 
                           X_Logic0_port, d(70) => X_Logic0_port, d(69) => 
                           X_Logic0_port, d(68) => X_Logic0_port, d(67) => 
                           X_Logic0_port, d(66) => X_Logic0_port, d(65) => 
                           X_Logic0_port, d(64) => X_Logic0_port, d(63) => 
                           X_Logic0_port, d(62) => X_Logic0_port, d(61) => 
                           X_Logic0_port, d(60) => X_Logic0_port, d(59) => 
                           X_Logic0_port, d(58) => X_Logic0_port, d(57) => 
                           X_Logic0_port, d(56) => X_Logic0_port, d(55) => 
                           X_Logic0_port, d(54) => X_Logic0_port, d(53) => 
                           X_Logic0_port, d(52) => X_Logic0_port, d(51) => 
                           X_Logic0_port, d(50) => X_Logic0_port, d(49) => 
                           X_Logic0_port, d(48) => X_Logic0_port, d(47) => 
                           X_Logic0_port, d(46) => X_Logic0_port, d(45) => 
                           X_Logic0_port, d(44) => X_Logic0_port, d(43) => 
                           X_Logic0_port, d(42) => X_Logic0_port, d(41) => 
                           X_Logic0_port, d(40) => X_Logic0_port, d(39) => 
                           X_Logic0_port, d(38) => X_Logic0_port, d(37) => 
                           X_Logic0_port, d(36) => X_Logic0_port, d(35) => 
                           X_Logic0_port, d(34) => X_Logic0_port, d(33) => 
                           X_Logic0_port, d(32) => X_Logic0_port, d(31) => 
                           X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           X_Logic0_port, d(20) => X_Logic0_port, d(19) => 
                           X_Logic0_port, d(18) => X_Logic0_port, d(17) => 
                           X_Logic0_port, d(16) => X_Logic0_port, d(15) => 
                           X_Logic0_port, d(14) => X_Logic0_port, d(13) => 
                           X_Logic0_port, d(12) => X_Logic0_port, d(11) => 
                           X_Logic0_port, d(10) => X_Logic0_port, d(9) => 
                           X_Logic0_port, d(8) => X_Logic0_port, d(7) => 
                           X_Logic0_port, d(6) => X_Logic0_port, d(5) => 
                           X_Logic0_port, d(4) => X_Logic0_port, d(3) => 
                           X_Logic0_port, d(2) => X_Logic0_port, d(1) => 
                           X_Logic0_port, d(0) => X_Logic0_port, Q(248) => 
                           n_3370, Q(247) => n_3371, Q(246) => n_3372, Q(245) 
                           => n_3373, Q(244) => n_3374, Q(243) => n_3375, 
                           Q(242) => n_3376, Q(241) => n_3377, Q(240) => n_3378
                           , Q(239) => n_3379, Q(238) => n_3380, Q(237) => 
                           n_3381, Q(236) => n_3382, Q(235) => n_3383, Q(234) 
                           => n_3384, Q(233) => n_3385, Q(232) => n_3386, 
                           Q(231) => n_3387, Q(230) => n_3388, Q(229) => n_3389
                           , Q(228) => n_3390, Q(227) => muxes_in_3_23_port, 
                           Q(226) => muxes_in_3_24_port, Q(225) => 
                           muxes_in_3_25_port, Q(224) => muxes_in_3_26_port, 
                           Q(223) => muxes_in_3_27_port, Q(222) => 
                           muxes_in_3_28_port, Q(221) => muxes_in_3_29_port, 
                           Q(220) => muxes_in_3_30_port, Q(219) => 
                           muxes_in_3_31_port, Q(218) => muxes_in_3_32_port, 
                           Q(217) => muxes_in_3_33_port, Q(216) => 
                           muxes_in_3_34_port, Q(215) => muxes_in_3_35_port, 
                           Q(214) => muxes_in_3_36_port, Q(213) => 
                           muxes_in_3_37_port, Q(212) => muxes_in_3_38_port, 
                           Q(211) => muxes_in_3_39_port, Q(210) => 
                           muxes_in_3_40_port, Q(209) => muxes_in_3_41_port, 
                           Q(208) => muxes_in_3_42_port, Q(207) => 
                           muxes_in_3_43_port, Q(206) => muxes_in_3_46_port, 
                           Q(205) => muxes_in_3_47_port, Q(204) => 
                           muxes_in_3_48_port, Q(203) => muxes_in_3_49_port, 
                           Q(202) => muxes_in_3_50_port, Q(201) => 
                           muxes_in_3_51_port, Q(200) => muxes_in_3_52_port, 
                           Q(199) => muxes_in_3_53_port, Q(198) => 
                           muxes_in_3_54_port, Q(197) => muxes_in_3_55_port, 
                           Q(196) => muxes_in_3_56_port, Q(195) => 
                           muxes_in_3_57_port, Q(194) => muxes_in_3_58_port, 
                           Q(193) => muxes_in_3_59_port, Q(192) => 
                           muxes_in_3_60_port, Q(191) => muxes_in_3_61_port, 
                           Q(190) => muxes_in_3_62_port, Q(189) => 
                           muxes_in_3_63_port, Q(188) => muxes_in_3_64_port, 
                           Q(187) => muxes_in_3_65_port, Q(186) => 
                           muxes_in_3_66_port, Q(185) => n_3391, Q(184) => 
                           n_3392, Q(183) => n_3393, Q(182) => n_3394, Q(181) 
                           => n_3395, Q(180) => n_3396, Q(179) => n_3397, 
                           Q(178) => n_3398, Q(177) => n_3399, Q(176) => n_3400
                           , Q(175) => n_3401, Q(174) => n_3402, Q(173) => 
                           n_3403, Q(172) => n_3404, Q(171) => n_3405, Q(170) 
                           => n_3406, Q(169) => n_3407, Q(168) => n_3408, 
                           Q(167) => n_3409, Q(166) => n_3410, Q(165) => n_3411
                           , Q(164) => n_3412, Q(163) => n_3413, Q(162) => 
                           n_3414, Q(161) => n_3415, Q(160) => n_3416, Q(159) 
                           => n_3417, Q(158) => n_3418, Q(157) => n_3419, 
                           Q(156) => n_3420, Q(155) => n_3421, Q(154) => n_3422
                           , Q(153) => n_3423, Q(152) => n_3424, Q(151) => 
                           n_3425, Q(150) => n_3426, Q(149) => n_3427, Q(148) 
                           => n_3428, Q(147) => n_3429, Q(146) => n_3430, 
                           Q(145) => n_3431, Q(144) => n_3432, Q(143) => n_3433
                           , Q(142) => n_3434, Q(141) => n_3435, Q(140) => 
                           n_3436, Q(139) => n_3437, Q(138) => n_3438, Q(137) 
                           => n_3439, Q(136) => n_3440, Q(135) => n_3441, 
                           Q(134) => n_3442, Q(133) => n_3443, Q(132) => n_3444
                           , Q(131) => n_3445, Q(130) => n_3446, Q(129) => 
                           n_3447, Q(128) => n_3448, Q(127) => n_3449, Q(126) 
                           => n_3450, Q(125) => n_3451, Q(124) => n_3452, 
                           Q(123) => n_3453, Q(122) => muxes_in_3_138_port, 
                           Q(121) => muxes_in_3_139_port, Q(120) => 
                           muxes_in_3_140_port, Q(119) => muxes_in_3_141_port, 
                           Q(118) => muxes_in_3_142_port, Q(117) => 
                           muxes_in_3_143_port, Q(116) => muxes_in_3_144_port, 
                           Q(115) => muxes_in_3_145_port, Q(114) => 
                           muxes_in_3_146_port, Q(113) => muxes_in_3_147_port, 
                           Q(112) => muxes_in_3_148_port, Q(111) => 
                           muxes_in_3_149_port, Q(110) => muxes_in_3_150_port, 
                           Q(109) => muxes_in_3_151_port, Q(108) => 
                           muxes_in_3_152_port, Q(107) => muxes_in_3_153_port, 
                           Q(106) => muxes_in_3_154_port, Q(105) => 
                           muxes_in_3_155_port, Q(104) => muxes_in_3_156_port, 
                           Q(103) => muxes_in_3_157_port, Q(102) => 
                           muxes_in_3_158_port, Q(101) => muxes_in_3_161_port, 
                           Q(100) => muxes_in_3_162_port, Q(99) => 
                           muxes_in_3_163_port, Q(98) => muxes_in_3_164_port, 
                           Q(97) => muxes_in_3_165_port, Q(96) => 
                           muxes_in_3_166_port, Q(95) => muxes_in_3_167_port, 
                           Q(94) => muxes_in_3_168_port, Q(93) => 
                           muxes_in_3_169_port, Q(92) => muxes_in_3_170_port, 
                           Q(91) => muxes_in_3_171_port, Q(90) => 
                           muxes_in_3_172_port, Q(89) => muxes_in_3_173_port, 
                           Q(88) => muxes_in_3_174_port, Q(87) => 
                           muxes_in_3_175_port, Q(86) => muxes_in_3_176_port, 
                           Q(85) => muxes_in_3_177_port, Q(84) => 
                           muxes_in_3_178_port, Q(83) => muxes_in_3_179_port, 
                           Q(82) => muxes_in_3_180_port, Q(81) => 
                           muxes_in_3_181_port, Q(80) => n_3454, Q(79) => 
                           n_3455, Q(78) => n_3456, Q(77) => n_3457, Q(76) => 
                           n_3458, Q(75) => n_3459, Q(74) => n_3460, Q(73) => 
                           n_3461, Q(72) => n_3462, Q(71) => n_3463, Q(70) => 
                           n_3464, Q(69) => n_3465, Q(68) => n_3466, Q(67) => 
                           n_3467, Q(66) => n_3468, Q(65) => n_3469, Q(64) => 
                           n_3470, Q(63) => n_3471, Q(62) => n_3472, Q(61) => 
                           n_3473, Q(60) => n_3474, Q(59) => n_3475, Q(58) => 
                           n_3476, Q(57) => n_3477, Q(56) => n_3478, Q(55) => 
                           n_3479, Q(54) => n_3480, Q(53) => n_3481, Q(52) => 
                           n_3482, Q(51) => n_3483, Q(50) => n_3484, Q(49) => 
                           n_3485, Q(48) => n_3486, Q(47) => n_3487, Q(46) => 
                           n_3488, Q(45) => n_3489, Q(44) => n_3490, Q(43) => 
                           n_3491, Q(42) => n_3492, Q(41) => n_3493, Q(40) => 
                           n_3494, Q(39) => n_3495, Q(38) => n_3496, Q(37) => 
                           n_3497, Q(36) => n_3498, Q(35) => n_3499, Q(34) => 
                           n_3500, Q(33) => n_3501, Q(32) => n_3502, Q(31) => 
                           n_3503, Q(30) => n_3504, Q(29) => n_3505, Q(28) => 
                           n_3506, Q(27) => n_3507, Q(26) => n_3508, Q(25) => 
                           n_3509, Q(24) => n_3510, Q(23) => n_3511, Q(22) => 
                           n_3512, Q(21) => n_3513, Q(20) => n_3514, Q(19) => 
                           n_3515, Q(18) => n_3516, Q(17) => n_3517, Q(16) => 
                           n_3518, Q(15) => n_3519, Q(14) => n_3520, Q(13) => 
                           n_3521, Q(12) => n_3522, Q(11) => n_3523, Q(10) => 
                           n_3524, Q(9) => n_3525, Q(8) => n_3526, Q(7) => 
                           n_3527, Q(6) => n_3528, Q(5) => n_3529, Q(4) => 
                           n_3530, Q(3) => n_3531, Q(2) => n_3532, Q(1) => 
                           n_3533, Q(0) => n_3534);
   MUXi_2 : MUX_zbit_nbit_N21_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           multiplier(15), inputs(22) => multiplier(15), 
                           inputs(23) => multiplier(14), inputs(24) => 
                           multiplier(13), inputs(25) => multiplier(12), 
                           inputs(26) => multiplier(11), inputs(27) => 
                           multiplier(10), inputs(28) => multiplier(9), 
                           inputs(29) => multiplier(8), inputs(30) => 
                           multiplier(7), inputs(31) => multiplier(6), 
                           inputs(32) => multiplier(5), inputs(33) => 
                           multiplier(4), inputs(34) => multiplier(3), 
                           inputs(35) => multiplier(2), inputs(36) => 
                           multiplier(1), inputs(37) => multiplier(0), 
                           inputs(38) => X_Logic0_port, inputs(39) => 
                           X_Logic0_port, inputs(40) => X_Logic0_port, 
                           inputs(41) => X_Logic0_port, inputs(42) => 
                           multiplier(15), inputs(43) => multiplier(14), 
                           inputs(44) => multiplier(13), inputs(45) => 
                           multiplier(12), inputs(46) => multiplier(11), 
                           inputs(47) => multiplier(10), inputs(48) => 
                           multiplier(9), inputs(49) => multiplier(8), 
                           inputs(50) => multiplier(7), inputs(51) => 
                           multiplier(6), inputs(52) => multiplier(5), 
                           inputs(53) => multiplier(4), inputs(54) => 
                           multiplier(3), inputs(55) => multiplier(2), 
                           inputs(56) => multiplier(1), inputs(57) => 
                           multiplier(0), inputs(58) => X_Logic0_port, 
                           inputs(59) => X_Logic0_port, inputs(60) => 
                           X_Logic0_port, inputs(61) => X_Logic0_port, 
                           inputs(62) => X_Logic0_port, inputs(63) => 
                           X_Logic0_port, inputs(64) => X_Logic0_port, 
                           inputs(65) => X_Logic0_port, inputs(66) => 
                           X_Logic0_port, inputs(67) => X_Logic0_port, 
                           inputs(68) => X_Logic0_port, inputs(69) => 
                           X_Logic0_port, inputs(70) => X_Logic0_port, 
                           inputs(71) => X_Logic0_port, inputs(72) => 
                           X_Logic0_port, inputs(73) => X_Logic0_port, 
                           inputs(74) => X_Logic0_port, inputs(75) => 
                           X_Logic0_port, inputs(76) => X_Logic0_port, 
                           inputs(77) => X_Logic0_port, inputs(78) => 
                           X_Logic0_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           muxes_in_0_102_port, inputs(127) => 
                           muxes_in_0_103_port, inputs(128) => 
                           muxes_in_0_104_port, inputs(129) => 
                           muxes_in_0_105_port, inputs(130) => 
                           muxes_in_0_106_port, inputs(131) => 
                           muxes_in_0_107_port, inputs(132) => 
                           muxes_in_0_108_port, inputs(133) => 
                           muxes_in_0_109_port, inputs(134) => 
                           muxes_in_0_110_port, inputs(135) => 
                           muxes_in_0_111_port, inputs(136) => 
                           muxes_in_0_112_port, inputs(137) => 
                           muxes_in_0_113_port, inputs(138) => 
                           muxes_in_0_114_port, inputs(139) => 
                           muxes_in_0_115_port, inputs(140) => 
                           muxes_in_0_116_port, inputs(141) => 
                           muxes_in_0_117_port, inputs(142) => X_Logic0_port, 
                           inputs(143) => X_Logic0_port, inputs(144) => 
                           X_Logic0_port, inputs(145) => X_Logic0_port, 
                           inputs(146) => X_Logic0_port, inputs(147) => 
                           muxes_in_0_119_port, inputs(148) => 
                           muxes_in_0_102_port, inputs(149) => 
                           muxes_in_0_103_port, inputs(150) => 
                           muxes_in_0_104_port, inputs(151) => 
                           muxes_in_0_105_port, inputs(152) => 
                           muxes_in_0_106_port, inputs(153) => 
                           muxes_in_0_107_port, inputs(154) => 
                           muxes_in_0_108_port, inputs(155) => 
                           muxes_in_0_109_port, inputs(156) => 
                           muxes_in_0_110_port, inputs(157) => 
                           muxes_in_0_111_port, inputs(158) => 
                           muxes_in_0_112_port, inputs(159) => 
                           muxes_in_0_113_port, inputs(160) => 
                           muxes_in_0_114_port, inputs(161) => 
                           muxes_in_0_115_port, inputs(162) => 
                           muxes_in_0_116_port, inputs(163) => 
                           muxes_in_0_117_port, inputs(164) => X_Logic0_port, 
                           inputs(165) => X_Logic0_port, inputs(166) => 
                           X_Logic0_port, inputs(167) => X_Logic0_port, SEL(2) 
                           => encoder_out_2_2_port, SEL(1) => 
                           encoder_out_2_1_port, SEL(0) => encoder_out_2_0_port
                           , Y(20) => mux_out_2_20_port, Y(19) => 
                           mux_out_2_19_port, Y(18) => mux_out_2_18_port, Y(17)
                           => mux_out_2_17_port, Y(16) => mux_out_2_16_port, 
                           Y(15) => mux_out_2_15_port, Y(14) => 
                           mux_out_2_14_port, Y(13) => mux_out_2_13_port, Y(12)
                           => mux_out_2_12_port, Y(11) => mux_out_2_11_port, 
                           Y(10) => mux_out_2_10_port, Y(9) => mux_out_2_9_port
                           , Y(8) => mux_out_2_8_port, Y(7) => mux_out_2_7_port
                           , Y(6) => mux_out_2_6_port, Y(5) => mux_out_2_5_port
                           , Y(4) => mux_out_2_4_port, Y(3) => mux_out_2_3_port
                           , Y(2) => mux_out_2_2_port, Y(1) => mux_out_2_1_port
                           , Y(0) => mux_out_2_0_port);
   ADDi_2 : adder_NBIT21 port map( a(20) => mux_out_2_20_port, a(19) => 
                           mux_out_2_19_port, a(18) => mux_out_2_18_port, a(17)
                           => mux_out_2_17_port, a(16) => mux_out_2_16_port, 
                           a(15) => mux_out_2_15_port, a(14) => 
                           mux_out_2_14_port, a(13) => mux_out_2_13_port, a(12)
                           => mux_out_2_12_port, a(11) => mux_out_2_11_port, 
                           a(10) => mux_out_2_10_port, a(9) => mux_out_2_9_port
                           , a(8) => mux_out_2_8_port, a(7) => mux_out_2_7_port
                           , a(6) => mux_out_2_6_port, a(5) => mux_out_2_5_port
                           , a(4) => mux_out_2_4_port, a(3) => mux_out_2_3_port
                           , a(2) => mux_out_2_2_port, a(1) => mux_out_2_1_port
                           , a(0) => mux_out_2_0_port, b(20) => 
                           sum_B_in_2_20_port, b(19) => sum_B_in_2_20_port, 
                           b(18) => sum_B_in_2_20_port, b(17) => 
                           sum_B_in_2_17_port, b(16) => sum_B_in_2_16_port, 
                           b(15) => sum_B_in_2_15_port, b(14) => 
                           sum_B_in_2_14_port, b(13) => sum_B_in_2_13_port, 
                           b(12) => sum_B_in_2_12_port, b(11) => 
                           sum_B_in_2_11_port, b(10) => sum_B_in_2_10_port, 
                           b(9) => sum_B_in_2_9_port, b(8) => sum_B_in_2_8_port
                           , b(7) => sum_B_in_2_7_port, b(6) => 
                           sum_B_in_2_6_port, b(5) => sum_B_in_2_5_port, b(4) 
                           => sum_B_in_2_4_port, b(3) => sum_B_in_2_3_port, 
                           b(2) => sum_B_in_2_2_port, b(1) => sum_B_in_2_1_port
                           , b(0) => sum_B_in_2_0_port, cin => X_Logic0_port, 
                           s(21) => sum_out_2_21_port, s(20) => 
                           sum_out_2_20_port, s(19) => sum_out_2_19_port, s(18)
                           => sum_out_2_18_port, s(17) => sum_out_2_17_port, 
                           s(16) => sum_out_2_16_port, s(15) => 
                           sum_out_2_15_port, s(14) => sum_out_2_14_port, s(13)
                           => sum_out_2_13_port, s(12) => sum_out_2_12_port, 
                           s(11) => sum_out_2_11_port, s(10) => 
                           sum_out_2_10_port, s(9) => sum_out_2_9_port, s(8) =>
                           sum_out_2_8_port, s(7) => sum_out_2_7_port, s(6) => 
                           sum_out_2_6_port, s(5) => sum_out_2_5_port, s(4) => 
                           sum_out_2_4_port, s(3) => sum_out_2_3_port, s(2) => 
                           sum_out_2_2_port, s(1) => sum_out_2_1_port, s(0) => 
                           sum_out_2_0_port);
   pip_del_reg_addi_2 : reg_nbit_n32_5 port map( clk => n12, reset => n5, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           sum_out_2_21_port, d(20) => sum_out_2_20_port, d(19)
                           => sum_out_2_19_port, d(18) => sum_out_2_18_port, 
                           d(17) => sum_out_2_17_port, d(16) => 
                           sum_out_2_16_port, d(15) => sum_out_2_15_port, d(14)
                           => sum_out_2_14_port, d(13) => sum_out_2_13_port, 
                           d(12) => sum_out_2_12_port, d(11) => 
                           sum_out_2_11_port, d(10) => sum_out_2_10_port, d(9) 
                           => sum_out_2_9_port, d(8) => sum_out_2_8_port, d(7) 
                           => sum_out_2_7_port, d(6) => sum_out_2_6_port, d(5) 
                           => sum_out_2_5_port, d(4) => sum_out_2_4_port, d(3) 
                           => sum_out_2_3_port, d(2) => sum_out_2_2_port, d(1) 
                           => sum_out_2_1_port, d(0) => sum_out_2_0_port, Q(31)
                           => n_3535, Q(30) => n_3536, Q(29) => n_3537, Q(28) 
                           => n_3538, Q(27) => n_3539, Q(26) => n_3540, Q(25) 
                           => n_3541, Q(24) => n_3542, Q(23) => n_3543, Q(22) 
                           => n_3544, Q(21) => n_3545, Q(20) => 
                           sum_B_in_3_22_port, Q(19) => sum_B_in_3_19_port, 
                           Q(18) => sum_B_in_3_18_port, Q(17) => 
                           sum_B_in_3_17_port, Q(16) => sum_B_in_3_16_port, 
                           Q(15) => sum_B_in_3_15_port, Q(14) => 
                           sum_B_in_3_14_port, Q(13) => sum_B_in_3_13_port, 
                           Q(12) => sum_B_in_3_12_port, Q(11) => 
                           sum_B_in_3_11_port, Q(10) => sum_B_in_3_10_port, 
                           Q(9) => sum_B_in_3_9_port, Q(8) => sum_B_in_3_8_port
                           , Q(7) => sum_B_in_3_7_port, Q(6) => 
                           sum_B_in_3_6_port, Q(5) => sum_B_in_3_5_port, Q(4) 
                           => sum_B_in_3_4_port, Q(3) => sum_B_in_3_3_port, 
                           Q(2) => sum_B_in_3_2_port, Q(1) => sum_B_in_3_1_port
                           , Q(0) => sum_B_in_3_0_port);
   ENCi_3 : encoder_5 port map( y(2) => multiplicand_pip_3_7_port, y(1) => 
                           multiplicand_pip_3_6_port, y(0) => 
                           multiplicand_pip_3_5_port, sel(2) => 
                           encoder_out_3_2_port, sel(1) => encoder_out_3_1_port
                           , sel(0) => encoder_out_3_0_port);
   pip_del_reg_muxi_3 : reg_nbit_n249_5 port map( clk => n10, reset => n5, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => X_Logic0_port, 
                           d(226) => X_Logic0_port, d(225) => 
                           muxes_in_3_23_port, d(224) => muxes_in_3_24_port, 
                           d(223) => muxes_in_3_25_port, d(222) => 
                           muxes_in_3_26_port, d(221) => muxes_in_3_27_port, 
                           d(220) => muxes_in_3_28_port, d(219) => 
                           muxes_in_3_29_port, d(218) => muxes_in_3_30_port, 
                           d(217) => muxes_in_3_31_port, d(216) => 
                           muxes_in_3_32_port, d(215) => muxes_in_3_33_port, 
                           d(214) => muxes_in_3_34_port, d(213) => 
                           muxes_in_3_35_port, d(212) => muxes_in_3_36_port, 
                           d(211) => muxes_in_3_37_port, d(210) => 
                           muxes_in_3_38_port, d(209) => muxes_in_3_39_port, 
                           d(208) => muxes_in_3_40_port, d(207) => 
                           muxes_in_3_41_port, d(206) => muxes_in_3_42_port, 
                           d(205) => muxes_in_3_43_port, d(204) => 
                           X_Logic0_port, d(203) => X_Logic0_port, d(202) => 
                           muxes_in_3_46_port, d(201) => muxes_in_3_47_port, 
                           d(200) => muxes_in_3_48_port, d(199) => 
                           muxes_in_3_49_port, d(198) => muxes_in_3_50_port, 
                           d(197) => muxes_in_3_51_port, d(196) => 
                           muxes_in_3_52_port, d(195) => muxes_in_3_53_port, 
                           d(194) => muxes_in_3_54_port, d(193) => 
                           muxes_in_3_55_port, d(192) => muxes_in_3_56_port, 
                           d(191) => muxes_in_3_57_port, d(190) => 
                           muxes_in_3_58_port, d(189) => muxes_in_3_59_port, 
                           d(188) => muxes_in_3_60_port, d(187) => 
                           muxes_in_3_61_port, d(186) => muxes_in_3_62_port, 
                           d(185) => muxes_in_3_63_port, d(184) => 
                           muxes_in_3_64_port, d(183) => muxes_in_3_65_port, 
                           d(182) => muxes_in_3_66_port, d(181) => 
                           X_Logic0_port, d(180) => X_Logic0_port, d(179) => 
                           X_Logic0_port, d(178) => X_Logic0_port, d(177) => 
                           X_Logic0_port, d(176) => X_Logic0_port, d(175) => 
                           X_Logic0_port, d(174) => X_Logic0_port, d(173) => 
                           X_Logic0_port, d(172) => X_Logic0_port, d(171) => 
                           X_Logic0_port, d(170) => X_Logic0_port, d(169) => 
                           X_Logic0_port, d(168) => X_Logic0_port, d(167) => 
                           X_Logic0_port, d(166) => X_Logic0_port, d(165) => 
                           X_Logic0_port, d(164) => X_Logic0_port, d(163) => 
                           X_Logic0_port, d(162) => X_Logic0_port, d(161) => 
                           X_Logic0_port, d(160) => X_Logic0_port, d(159) => 
                           X_Logic0_port, d(158) => X_Logic0_port, d(157) => 
                           X_Logic0_port, d(156) => X_Logic0_port, d(155) => 
                           X_Logic0_port, d(154) => X_Logic0_port, d(153) => 
                           X_Logic0_port, d(152) => X_Logic0_port, d(151) => 
                           X_Logic0_port, d(150) => X_Logic0_port, d(149) => 
                           X_Logic0_port, d(148) => X_Logic0_port, d(147) => 
                           X_Logic0_port, d(146) => X_Logic0_port, d(145) => 
                           X_Logic0_port, d(144) => X_Logic0_port, d(143) => 
                           X_Logic0_port, d(142) => X_Logic0_port, d(141) => 
                           X_Logic0_port, d(140) => X_Logic0_port, d(139) => 
                           X_Logic0_port, d(138) => X_Logic0_port, d(137) => 
                           X_Logic0_port, d(136) => X_Logic0_port, d(135) => 
                           X_Logic0_port, d(134) => X_Logic0_port, d(133) => 
                           X_Logic0_port, d(132) => X_Logic0_port, d(131) => 
                           X_Logic0_port, d(130) => X_Logic0_port, d(129) => 
                           X_Logic0_port, d(128) => X_Logic0_port, d(127) => 
                           X_Logic0_port, d(126) => X_Logic0_port, d(125) => 
                           X_Logic0_port, d(124) => X_Logic0_port, d(123) => 
                           X_Logic0_port, d(122) => X_Logic0_port, d(121) => 
                           X_Logic0_port, d(120) => X_Logic0_port, d(119) => 
                           X_Logic0_port, d(118) => X_Logic0_port, d(117) => 
                           X_Logic0_port, d(116) => X_Logic0_port, d(115) => 
                           X_Logic0_port, d(114) => X_Logic0_port, d(113) => 
                           X_Logic0_port, d(112) => X_Logic0_port, d(111) => 
                           X_Logic0_port, d(110) => muxes_in_3_138_port, d(109)
                           => muxes_in_3_139_port, d(108) => 
                           muxes_in_3_140_port, d(107) => muxes_in_3_141_port, 
                           d(106) => muxes_in_3_142_port, d(105) => 
                           muxes_in_3_143_port, d(104) => muxes_in_3_144_port, 
                           d(103) => muxes_in_3_145_port, d(102) => 
                           muxes_in_3_146_port, d(101) => muxes_in_3_147_port, 
                           d(100) => muxes_in_3_148_port, d(99) => 
                           muxes_in_3_149_port, d(98) => muxes_in_3_150_port, 
                           d(97) => muxes_in_3_151_port, d(96) => 
                           muxes_in_3_152_port, d(95) => muxes_in_3_153_port, 
                           d(94) => muxes_in_3_154_port, d(93) => 
                           muxes_in_3_155_port, d(92) => muxes_in_3_156_port, 
                           d(91) => muxes_in_3_157_port, d(90) => 
                           muxes_in_3_158_port, d(89) => X_Logic0_port, d(88) 
                           => X_Logic0_port, d(87) => muxes_in_3_161_port, 
                           d(86) => muxes_in_3_162_port, d(85) => 
                           muxes_in_3_163_port, d(84) => muxes_in_3_164_port, 
                           d(83) => muxes_in_3_165_port, d(82) => 
                           muxes_in_3_166_port, d(81) => muxes_in_3_167_port, 
                           d(80) => muxes_in_3_168_port, d(79) => 
                           muxes_in_3_169_port, d(78) => muxes_in_3_170_port, 
                           d(77) => muxes_in_3_171_port, d(76) => 
                           muxes_in_3_172_port, d(75) => muxes_in_3_173_port, 
                           d(74) => muxes_in_3_174_port, d(73) => 
                           muxes_in_3_175_port, d(72) => muxes_in_3_176_port, 
                           d(71) => muxes_in_3_177_port, d(70) => 
                           muxes_in_3_178_port, d(69) => muxes_in_3_179_port, 
                           d(68) => muxes_in_3_180_port, d(67) => 
                           muxes_in_3_181_port, d(66) => X_Logic0_port, d(65) 
                           => X_Logic0_port, d(64) => X_Logic0_port, d(63) => 
                           X_Logic0_port, d(62) => X_Logic0_port, d(61) => 
                           X_Logic0_port, d(60) => X_Logic0_port, d(59) => 
                           X_Logic0_port, d(58) => X_Logic0_port, d(57) => 
                           X_Logic0_port, d(56) => X_Logic0_port, d(55) => 
                           X_Logic0_port, d(54) => X_Logic0_port, d(53) => 
                           X_Logic0_port, d(52) => X_Logic0_port, d(51) => 
                           X_Logic0_port, d(50) => X_Logic0_port, d(49) => 
                           X_Logic0_port, d(48) => X_Logic0_port, d(47) => 
                           X_Logic0_port, d(46) => X_Logic0_port, d(45) => 
                           X_Logic0_port, d(44) => X_Logic0_port, d(43) => 
                           X_Logic0_port, d(42) => X_Logic0_port, d(41) => 
                           X_Logic0_port, d(40) => X_Logic0_port, d(39) => 
                           X_Logic0_port, d(38) => X_Logic0_port, d(37) => 
                           X_Logic0_port, d(36) => X_Logic0_port, d(35) => 
                           X_Logic0_port, d(34) => X_Logic0_port, d(33) => 
                           X_Logic0_port, d(32) => X_Logic0_port, d(31) => 
                           X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           X_Logic0_port, d(20) => X_Logic0_port, d(19) => 
                           X_Logic0_port, d(18) => X_Logic0_port, d(17) => 
                           X_Logic0_port, d(16) => X_Logic0_port, d(15) => 
                           X_Logic0_port, d(14) => X_Logic0_port, d(13) => 
                           X_Logic0_port, d(12) => X_Logic0_port, d(11) => 
                           X_Logic0_port, d(10) => X_Logic0_port, d(9) => 
                           X_Logic0_port, d(8) => X_Logic0_port, d(7) => 
                           X_Logic0_port, d(6) => X_Logic0_port, d(5) => 
                           X_Logic0_port, d(4) => X_Logic0_port, d(3) => 
                           X_Logic0_port, d(2) => X_Logic0_port, d(1) => 
                           X_Logic0_port, d(0) => X_Logic0_port, Q(248) => 
                           n_3546, Q(247) => n_3547, Q(246) => n_3548, Q(245) 
                           => n_3549, Q(244) => n_3550, Q(243) => n_3551, 
                           Q(242) => n_3552, Q(241) => n_3553, Q(240) => n_3554
                           , Q(239) => n_3555, Q(238) => n_3556, Q(237) => 
                           n_3557, Q(236) => n_3558, Q(235) => n_3559, Q(234) 
                           => n_3560, Q(233) => n_3561, Q(232) => n_3562, 
                           Q(231) => n_3563, Q(230) => n_3564, Q(229) => n_3565
                           , Q(228) => n_3566, Q(227) => n_3567, Q(226) => 
                           n_3568, Q(225) => muxes_in_4_25_port, Q(224) => 
                           muxes_in_4_26_port, Q(223) => muxes_in_4_27_port, 
                           Q(222) => muxes_in_4_28_port, Q(221) => 
                           muxes_in_4_29_port, Q(220) => muxes_in_4_30_port, 
                           Q(219) => muxes_in_4_31_port, Q(218) => 
                           muxes_in_4_32_port, Q(217) => muxes_in_4_33_port, 
                           Q(216) => muxes_in_4_34_port, Q(215) => 
                           muxes_in_4_35_port, Q(214) => muxes_in_4_36_port, 
                           Q(213) => muxes_in_4_37_port, Q(212) => 
                           muxes_in_4_38_port, Q(211) => muxes_in_4_39_port, 
                           Q(210) => muxes_in_4_40_port, Q(209) => 
                           muxes_in_4_41_port, Q(208) => muxes_in_4_42_port, 
                           Q(207) => muxes_in_4_43_port, Q(206) => 
                           muxes_in_4_44_port, Q(205) => muxes_in_4_45_port, 
                           Q(204) => muxes_in_4_46_port, Q(203) => 
                           muxes_in_4_47_port, Q(202) => muxes_in_4_50_port, 
                           Q(201) => muxes_in_4_51_port, Q(200) => 
                           muxes_in_4_52_port, Q(199) => muxes_in_4_53_port, 
                           Q(198) => muxes_in_4_54_port, Q(197) => 
                           muxes_in_4_55_port, Q(196) => muxes_in_4_56_port, 
                           Q(195) => muxes_in_4_57_port, Q(194) => 
                           muxes_in_4_58_port, Q(193) => muxes_in_4_59_port, 
                           Q(192) => muxes_in_4_60_port, Q(191) => 
                           muxes_in_4_61_port, Q(190) => muxes_in_4_62_port, 
                           Q(189) => muxes_in_4_63_port, Q(188) => 
                           muxes_in_4_64_port, Q(187) => muxes_in_4_65_port, 
                           Q(186) => muxes_in_4_66_port, Q(185) => 
                           muxes_in_4_67_port, Q(184) => muxes_in_4_68_port, 
                           Q(183) => muxes_in_4_69_port, Q(182) => 
                           muxes_in_4_70_port, Q(181) => muxes_in_4_71_port, 
                           Q(180) => muxes_in_4_72_port, Q(179) => n_3569, 
                           Q(178) => n_3570, Q(177) => n_3571, Q(176) => n_3572
                           , Q(175) => n_3573, Q(174) => n_3574, Q(173) => 
                           n_3575, Q(172) => n_3576, Q(171) => n_3577, Q(170) 
                           => n_3578, Q(169) => n_3579, Q(168) => n_3580, 
                           Q(167) => n_3581, Q(166) => n_3582, Q(165) => n_3583
                           , Q(164) => n_3584, Q(163) => n_3585, Q(162) => 
                           n_3586, Q(161) => n_3587, Q(160) => n_3588, Q(159) 
                           => n_3589, Q(158) => n_3590, Q(157) => n_3591, 
                           Q(156) => n_3592, Q(155) => n_3593, Q(154) => n_3594
                           , Q(153) => n_3595, Q(152) => n_3596, Q(151) => 
                           n_3597, Q(150) => n_3598, Q(149) => n_3599, Q(148) 
                           => n_3600, Q(147) => n_3601, Q(146) => n_3602, 
                           Q(145) => n_3603, Q(144) => n_3604, Q(143) => n_3605
                           , Q(142) => n_3606, Q(141) => n_3607, Q(140) => 
                           n_3608, Q(139) => n_3609, Q(138) => n_3610, Q(137) 
                           => n_3611, Q(136) => n_3612, Q(135) => n_3613, 
                           Q(134) => n_3614, Q(133) => n_3615, Q(132) => n_3616
                           , Q(131) => n_3617, Q(130) => n_3618, Q(129) => 
                           n_3619, Q(128) => n_3620, Q(127) => n_3621, Q(126) 
                           => n_3622, Q(125) => n_3623, Q(124) => n_3624, 
                           Q(123) => n_3625, Q(122) => n_3626, Q(121) => n_3627
                           , Q(120) => n_3628, Q(119) => n_3629, Q(118) => 
                           n_3630, Q(117) => n_3631, Q(116) => n_3632, Q(115) 
                           => n_3633, Q(114) => n_3634, Q(113) => n_3635, 
                           Q(112) => n_3636, Q(111) => n_3637, Q(110) => 
                           muxes_in_4_150_port, Q(109) => muxes_in_4_151_port, 
                           Q(108) => muxes_in_4_152_port, Q(107) => 
                           muxes_in_4_153_port, Q(106) => muxes_in_4_154_port, 
                           Q(105) => muxes_in_4_155_port, Q(104) => 
                           muxes_in_4_156_port, Q(103) => muxes_in_4_157_port, 
                           Q(102) => muxes_in_4_158_port, Q(101) => 
                           muxes_in_4_159_port, Q(100) => muxes_in_4_160_port, 
                           Q(99) => muxes_in_4_161_port, Q(98) => 
                           muxes_in_4_162_port, Q(97) => muxes_in_4_163_port, 
                           Q(96) => muxes_in_4_164_port, Q(95) => 
                           muxes_in_4_165_port, Q(94) => muxes_in_4_166_port, 
                           Q(93) => muxes_in_4_167_port, Q(92) => 
                           muxes_in_4_168_port, Q(91) => muxes_in_4_169_port, 
                           Q(90) => muxes_in_4_170_port, Q(89) => 
                           muxes_in_4_171_port, Q(88) => muxes_in_4_172_port, 
                           Q(87) => muxes_in_4_175_port, Q(86) => 
                           muxes_in_4_176_port, Q(85) => muxes_in_4_177_port, 
                           Q(84) => muxes_in_4_178_port, Q(83) => 
                           muxes_in_4_179_port, Q(82) => muxes_in_4_180_port, 
                           Q(81) => muxes_in_4_181_port, Q(80) => 
                           muxes_in_4_182_port, Q(79) => muxes_in_4_183_port, 
                           Q(78) => muxes_in_4_184_port, Q(77) => 
                           muxes_in_4_185_port, Q(76) => muxes_in_4_186_port, 
                           Q(75) => muxes_in_4_187_port, Q(74) => 
                           muxes_in_4_188_port, Q(73) => muxes_in_4_189_port, 
                           Q(72) => muxes_in_4_190_port, Q(71) => 
                           muxes_in_4_191_port, Q(70) => muxes_in_4_192_port, 
                           Q(69) => muxes_in_4_193_port, Q(68) => 
                           muxes_in_4_194_port, Q(67) => muxes_in_4_195_port, 
                           Q(66) => muxes_in_4_196_port, Q(65) => 
                           muxes_in_4_197_port, Q(64) => n_3638, Q(63) => 
                           n_3639, Q(62) => n_3640, Q(61) => n_3641, Q(60) => 
                           n_3642, Q(59) => n_3643, Q(58) => n_3644, Q(57) => 
                           n_3645, Q(56) => n_3646, Q(55) => n_3647, Q(54) => 
                           n_3648, Q(53) => n_3649, Q(52) => n_3650, Q(51) => 
                           n_3651, Q(50) => n_3652, Q(49) => n_3653, Q(48) => 
                           n_3654, Q(47) => n_3655, Q(46) => n_3656, Q(45) => 
                           n_3657, Q(44) => n_3658, Q(43) => n_3659, Q(42) => 
                           n_3660, Q(41) => n_3661, Q(40) => n_3662, Q(39) => 
                           n_3663, Q(38) => n_3664, Q(37) => n_3665, Q(36) => 
                           n_3666, Q(35) => n_3667, Q(34) => n_3668, Q(33) => 
                           n_3669, Q(32) => n_3670, Q(31) => n_3671, Q(30) => 
                           n_3672, Q(29) => n_3673, Q(28) => n_3674, Q(27) => 
                           n_3675, Q(26) => n_3676, Q(25) => n_3677, Q(24) => 
                           n_3678, Q(23) => n_3679, Q(22) => n_3680, Q(21) => 
                           n_3681, Q(20) => n_3682, Q(19) => n_3683, Q(18) => 
                           n_3684, Q(17) => n_3685, Q(16) => n_3686, Q(15) => 
                           n_3687, Q(14) => n_3688, Q(13) => n_3689, Q(12) => 
                           n_3690, Q(11) => n_3691, Q(10) => n_3692, Q(9) => 
                           n_3693, Q(8) => n_3694, Q(7) => n_3695, Q(6) => 
                           n_3696, Q(5) => n_3697, Q(4) => n_3698, Q(3) => 
                           n_3699, Q(2) => n_3700, Q(1) => n_3701, Q(0) => 
                           n_3702);
   MUXi_3 : MUX_zbit_nbit_N23_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           X_Logic0_port, inputs(22) => X_Logic0_port, 
                           inputs(23) => muxes_in_3_23_port, inputs(24) => 
                           muxes_in_3_24_port, inputs(25) => muxes_in_3_25_port
                           , inputs(26) => muxes_in_3_26_port, inputs(27) => 
                           muxes_in_3_27_port, inputs(28) => muxes_in_3_28_port
                           , inputs(29) => muxes_in_3_29_port, inputs(30) => 
                           muxes_in_3_30_port, inputs(31) => muxes_in_3_31_port
                           , inputs(32) => muxes_in_3_32_port, inputs(33) => 
                           muxes_in_3_33_port, inputs(34) => muxes_in_3_34_port
                           , inputs(35) => muxes_in_3_35_port, inputs(36) => 
                           muxes_in_3_36_port, inputs(37) => muxes_in_3_37_port
                           , inputs(38) => muxes_in_3_38_port, inputs(39) => 
                           muxes_in_3_39_port, inputs(40) => muxes_in_3_40_port
                           , inputs(41) => muxes_in_3_41_port, inputs(42) => 
                           muxes_in_3_42_port, inputs(43) => muxes_in_3_43_port
                           , inputs(44) => X_Logic0_port, inputs(45) => 
                           X_Logic0_port, inputs(46) => muxes_in_3_46_port, 
                           inputs(47) => muxes_in_3_47_port, inputs(48) => 
                           muxes_in_3_48_port, inputs(49) => muxes_in_3_49_port
                           , inputs(50) => muxes_in_3_50_port, inputs(51) => 
                           muxes_in_3_51_port, inputs(52) => muxes_in_3_52_port
                           , inputs(53) => muxes_in_3_53_port, inputs(54) => 
                           muxes_in_3_54_port, inputs(55) => muxes_in_3_55_port
                           , inputs(56) => muxes_in_3_56_port, inputs(57) => 
                           muxes_in_3_57_port, inputs(58) => muxes_in_3_58_port
                           , inputs(59) => muxes_in_3_59_port, inputs(60) => 
                           muxes_in_3_60_port, inputs(61) => muxes_in_3_61_port
                           , inputs(62) => muxes_in_3_62_port, inputs(63) => 
                           muxes_in_3_63_port, inputs(64) => muxes_in_3_64_port
                           , inputs(65) => muxes_in_3_65_port, inputs(66) => 
                           muxes_in_3_66_port, inputs(67) => X_Logic0_port, 
                           inputs(68) => X_Logic0_port, inputs(69) => 
                           X_Logic0_port, inputs(70) => X_Logic0_port, 
                           inputs(71) => X_Logic0_port, inputs(72) => 
                           X_Logic0_port, inputs(73) => X_Logic0_port, 
                           inputs(74) => X_Logic0_port, inputs(75) => 
                           X_Logic0_port, inputs(76) => X_Logic0_port, 
                           inputs(77) => X_Logic0_port, inputs(78) => 
                           X_Logic0_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           X_Logic0_port, inputs(127) => X_Logic0_port, 
                           inputs(128) => X_Logic0_port, inputs(129) => 
                           X_Logic0_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => X_Logic0_port, 
                           inputs(134) => X_Logic0_port, inputs(135) => 
                           X_Logic0_port, inputs(136) => X_Logic0_port, 
                           inputs(137) => X_Logic0_port, inputs(138) => 
                           muxes_in_3_138_port, inputs(139) => 
                           muxes_in_3_139_port, inputs(140) => 
                           muxes_in_3_140_port, inputs(141) => 
                           muxes_in_3_141_port, inputs(142) => 
                           muxes_in_3_142_port, inputs(143) => 
                           muxes_in_3_143_port, inputs(144) => 
                           muxes_in_3_144_port, inputs(145) => 
                           muxes_in_3_145_port, inputs(146) => 
                           muxes_in_3_146_port, inputs(147) => 
                           muxes_in_3_147_port, inputs(148) => 
                           muxes_in_3_148_port, inputs(149) => 
                           muxes_in_3_149_port, inputs(150) => 
                           muxes_in_3_150_port, inputs(151) => 
                           muxes_in_3_151_port, inputs(152) => 
                           muxes_in_3_152_port, inputs(153) => 
                           muxes_in_3_153_port, inputs(154) => 
                           muxes_in_3_154_port, inputs(155) => 
                           muxes_in_3_155_port, inputs(156) => 
                           muxes_in_3_156_port, inputs(157) => 
                           muxes_in_3_157_port, inputs(158) => 
                           muxes_in_3_158_port, inputs(159) => X_Logic0_port, 
                           inputs(160) => X_Logic0_port, inputs(161) => 
                           muxes_in_3_161_port, inputs(162) => 
                           muxes_in_3_162_port, inputs(163) => 
                           muxes_in_3_163_port, inputs(164) => 
                           muxes_in_3_164_port, inputs(165) => 
                           muxes_in_3_165_port, inputs(166) => 
                           muxes_in_3_166_port, inputs(167) => 
                           muxes_in_3_167_port, inputs(168) => 
                           muxes_in_3_168_port, inputs(169) => 
                           muxes_in_3_169_port, inputs(170) => 
                           muxes_in_3_170_port, inputs(171) => 
                           muxes_in_3_171_port, inputs(172) => 
                           muxes_in_3_172_port, inputs(173) => 
                           muxes_in_3_173_port, inputs(174) => 
                           muxes_in_3_174_port, inputs(175) => 
                           muxes_in_3_175_port, inputs(176) => 
                           muxes_in_3_176_port, inputs(177) => 
                           muxes_in_3_177_port, inputs(178) => 
                           muxes_in_3_178_port, inputs(179) => 
                           muxes_in_3_179_port, inputs(180) => 
                           muxes_in_3_180_port, inputs(181) => 
                           muxes_in_3_181_port, inputs(182) => X_Logic0_port, 
                           inputs(183) => X_Logic0_port, SEL(2) => 
                           encoder_out_3_2_port, SEL(1) => encoder_out_3_1_port
                           , SEL(0) => encoder_out_3_0_port, Y(22) => 
                           mux_out_3_22_port, Y(21) => mux_out_3_21_port, Y(20)
                           => mux_out_3_20_port, Y(19) => mux_out_3_19_port, 
                           Y(18) => mux_out_3_18_port, Y(17) => 
                           mux_out_3_17_port, Y(16) => mux_out_3_16_port, Y(15)
                           => mux_out_3_15_port, Y(14) => mux_out_3_14_port, 
                           Y(13) => mux_out_3_13_port, Y(12) => 
                           mux_out_3_12_port, Y(11) => mux_out_3_11_port, Y(10)
                           => mux_out_3_10_port, Y(9) => mux_out_3_9_port, Y(8)
                           => mux_out_3_8_port, Y(7) => mux_out_3_7_port, Y(6) 
                           => mux_out_3_6_port, Y(5) => mux_out_3_5_port, Y(4) 
                           => mux_out_3_4_port, Y(3) => mux_out_3_3_port, Y(2) 
                           => mux_out_3_2_port, Y(1) => mux_out_3_1_port, Y(0) 
                           => mux_out_3_0_port);
   ADDi_3 : adder_NBIT23 port map( a(22) => mux_out_3_22_port, a(21) => 
                           mux_out_3_21_port, a(20) => mux_out_3_20_port, a(19)
                           => mux_out_3_19_port, a(18) => mux_out_3_18_port, 
                           a(17) => mux_out_3_17_port, a(16) => 
                           mux_out_3_16_port, a(15) => mux_out_3_15_port, a(14)
                           => mux_out_3_14_port, a(13) => mux_out_3_13_port, 
                           a(12) => mux_out_3_12_port, a(11) => 
                           mux_out_3_11_port, a(10) => mux_out_3_10_port, a(9) 
                           => mux_out_3_9_port, a(8) => mux_out_3_8_port, a(7) 
                           => mux_out_3_7_port, a(6) => mux_out_3_6_port, a(5) 
                           => mux_out_3_5_port, a(4) => mux_out_3_4_port, a(3) 
                           => mux_out_3_3_port, a(2) => mux_out_3_2_port, a(1) 
                           => mux_out_3_1_port, a(0) => mux_out_3_0_port, b(22)
                           => sum_B_in_3_22_port, b(21) => sum_B_in_3_22_port, 
                           b(20) => sum_B_in_3_22_port, b(19) => 
                           sum_B_in_3_19_port, b(18) => sum_B_in_3_18_port, 
                           b(17) => sum_B_in_3_17_port, b(16) => 
                           sum_B_in_3_16_port, b(15) => sum_B_in_3_15_port, 
                           b(14) => sum_B_in_3_14_port, b(13) => 
                           sum_B_in_3_13_port, b(12) => sum_B_in_3_12_port, 
                           b(11) => sum_B_in_3_11_port, b(10) => 
                           sum_B_in_3_10_port, b(9) => sum_B_in_3_9_port, b(8) 
                           => sum_B_in_3_8_port, b(7) => sum_B_in_3_7_port, 
                           b(6) => sum_B_in_3_6_port, b(5) => sum_B_in_3_5_port
                           , b(4) => sum_B_in_3_4_port, b(3) => 
                           sum_B_in_3_3_port, b(2) => sum_B_in_3_2_port, b(1) 
                           => sum_B_in_3_1_port, b(0) => sum_B_in_3_0_port, cin
                           => X_Logic0_port, s(23) => sum_out_3_23_port, s(22) 
                           => sum_out_3_22_port, s(21) => sum_out_3_21_port, 
                           s(20) => sum_out_3_20_port, s(19) => 
                           sum_out_3_19_port, s(18) => sum_out_3_18_port, s(17)
                           => sum_out_3_17_port, s(16) => sum_out_3_16_port, 
                           s(15) => sum_out_3_15_port, s(14) => 
                           sum_out_3_14_port, s(13) => sum_out_3_13_port, s(12)
                           => sum_out_3_12_port, s(11) => sum_out_3_11_port, 
                           s(10) => sum_out_3_10_port, s(9) => sum_out_3_9_port
                           , s(8) => sum_out_3_8_port, s(7) => sum_out_3_7_port
                           , s(6) => sum_out_3_6_port, s(5) => sum_out_3_5_port
                           , s(4) => sum_out_3_4_port, s(3) => sum_out_3_3_port
                           , s(2) => sum_out_3_2_port, s(1) => sum_out_3_1_port
                           , s(0) => sum_out_3_0_port);
   pip_del_reg_addi_3 : reg_nbit_n32_4 port map( clk => n12, reset => n5, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           sum_out_3_23_port, d(22) => sum_out_3_22_port, d(21)
                           => sum_out_3_21_port, d(20) => sum_out_3_20_port, 
                           d(19) => sum_out_3_19_port, d(18) => 
                           sum_out_3_18_port, d(17) => sum_out_3_17_port, d(16)
                           => sum_out_3_16_port, d(15) => sum_out_3_15_port, 
                           d(14) => sum_out_3_14_port, d(13) => 
                           sum_out_3_13_port, d(12) => sum_out_3_12_port, d(11)
                           => sum_out_3_11_port, d(10) => sum_out_3_10_port, 
                           d(9) => sum_out_3_9_port, d(8) => sum_out_3_8_port, 
                           d(7) => sum_out_3_7_port, d(6) => sum_out_3_6_port, 
                           d(5) => sum_out_3_5_port, d(4) => sum_out_3_4_port, 
                           d(3) => sum_out_3_3_port, d(2) => sum_out_3_2_port, 
                           d(1) => sum_out_3_1_port, d(0) => sum_out_3_0_port, 
                           Q(31) => n_3703, Q(30) => n_3704, Q(29) => n_3705, 
                           Q(28) => n_3706, Q(27) => n_3707, Q(26) => n_3708, 
                           Q(25) => n_3709, Q(24) => n_3710, Q(23) => n_3711, 
                           Q(22) => sum_B_in_4_24_port, Q(21) => 
                           sum_B_in_4_21_port, Q(20) => sum_B_in_4_20_port, 
                           Q(19) => sum_B_in_4_19_port, Q(18) => 
                           sum_B_in_4_18_port, Q(17) => sum_B_in_4_17_port, 
                           Q(16) => sum_B_in_4_16_port, Q(15) => 
                           sum_B_in_4_15_port, Q(14) => sum_B_in_4_14_port, 
                           Q(13) => sum_B_in_4_13_port, Q(12) => 
                           sum_B_in_4_12_port, Q(11) => sum_B_in_4_11_port, 
                           Q(10) => sum_B_in_4_10_port, Q(9) => 
                           sum_B_in_4_9_port, Q(8) => sum_B_in_4_8_port, Q(7) 
                           => sum_B_in_4_7_port, Q(6) => sum_B_in_4_6_port, 
                           Q(5) => sum_B_in_4_5_port, Q(4) => sum_B_in_4_4_port
                           , Q(3) => sum_B_in_4_3_port, Q(2) => 
                           sum_B_in_4_2_port, Q(1) => sum_B_in_4_1_port, Q(0) 
                           => sum_B_in_4_0_port);
   ENCi_4 : encoder_4 port map( y(2) => multiplicand_pip_4_9_port, y(1) => 
                           multiplicand_pip_4_8_port, y(0) => 
                           multiplicand_pip_4_7_port, sel(2) => 
                           encoder_out_4_2_port, sel(1) => encoder_out_4_1_port
                           , sel(0) => encoder_out_4_0_port);
   pip_del_reg_muxi_4 : reg_nbit_n249_4 port map( clk => n10, reset => n5, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => X_Logic0_port, 
                           d(226) => X_Logic0_port, d(225) => X_Logic0_port, 
                           d(224) => X_Logic0_port, d(223) => 
                           muxes_in_4_25_port, d(222) => muxes_in_4_26_port, 
                           d(221) => muxes_in_4_27_port, d(220) => 
                           muxes_in_4_28_port, d(219) => muxes_in_4_29_port, 
                           d(218) => muxes_in_4_30_port, d(217) => 
                           muxes_in_4_31_port, d(216) => muxes_in_4_32_port, 
                           d(215) => muxes_in_4_33_port, d(214) => 
                           muxes_in_4_34_port, d(213) => muxes_in_4_35_port, 
                           d(212) => muxes_in_4_36_port, d(211) => 
                           muxes_in_4_37_port, d(210) => muxes_in_4_38_port, 
                           d(209) => muxes_in_4_39_port, d(208) => 
                           muxes_in_4_40_port, d(207) => muxes_in_4_41_port, 
                           d(206) => muxes_in_4_42_port, d(205) => 
                           muxes_in_4_43_port, d(204) => muxes_in_4_44_port, 
                           d(203) => muxes_in_4_45_port, d(202) => 
                           muxes_in_4_46_port, d(201) => muxes_in_4_47_port, 
                           d(200) => X_Logic0_port, d(199) => X_Logic0_port, 
                           d(198) => muxes_in_4_50_port, d(197) => 
                           muxes_in_4_51_port, d(196) => muxes_in_4_52_port, 
                           d(195) => muxes_in_4_53_port, d(194) => 
                           muxes_in_4_54_port, d(193) => muxes_in_4_55_port, 
                           d(192) => muxes_in_4_56_port, d(191) => 
                           muxes_in_4_57_port, d(190) => muxes_in_4_58_port, 
                           d(189) => muxes_in_4_59_port, d(188) => 
                           muxes_in_4_60_port, d(187) => muxes_in_4_61_port, 
                           d(186) => muxes_in_4_62_port, d(185) => 
                           muxes_in_4_63_port, d(184) => muxes_in_4_64_port, 
                           d(183) => muxes_in_4_65_port, d(182) => 
                           muxes_in_4_66_port, d(181) => muxes_in_4_67_port, 
                           d(180) => muxes_in_4_68_port, d(179) => 
                           muxes_in_4_69_port, d(178) => muxes_in_4_70_port, 
                           d(177) => muxes_in_4_71_port, d(176) => 
                           muxes_in_4_72_port, d(175) => X_Logic0_port, d(174) 
                           => X_Logic0_port, d(173) => X_Logic0_port, d(172) =>
                           X_Logic0_port, d(171) => X_Logic0_port, d(170) => 
                           X_Logic0_port, d(169) => X_Logic0_port, d(168) => 
                           X_Logic0_port, d(167) => X_Logic0_port, d(166) => 
                           X_Logic0_port, d(165) => X_Logic0_port, d(164) => 
                           X_Logic0_port, d(163) => X_Logic0_port, d(162) => 
                           X_Logic0_port, d(161) => X_Logic0_port, d(160) => 
                           X_Logic0_port, d(159) => X_Logic0_port, d(158) => 
                           X_Logic0_port, d(157) => X_Logic0_port, d(156) => 
                           X_Logic0_port, d(155) => X_Logic0_port, d(154) => 
                           X_Logic0_port, d(153) => X_Logic0_port, d(152) => 
                           X_Logic0_port, d(151) => X_Logic0_port, d(150) => 
                           X_Logic0_port, d(149) => X_Logic0_port, d(148) => 
                           X_Logic0_port, d(147) => X_Logic0_port, d(146) => 
                           X_Logic0_port, d(145) => X_Logic0_port, d(144) => 
                           X_Logic0_port, d(143) => X_Logic0_port, d(142) => 
                           X_Logic0_port, d(141) => X_Logic0_port, d(140) => 
                           X_Logic0_port, d(139) => X_Logic0_port, d(138) => 
                           X_Logic0_port, d(137) => X_Logic0_port, d(136) => 
                           X_Logic0_port, d(135) => X_Logic0_port, d(134) => 
                           X_Logic0_port, d(133) => X_Logic0_port, d(132) => 
                           X_Logic0_port, d(131) => X_Logic0_port, d(130) => 
                           X_Logic0_port, d(129) => X_Logic0_port, d(128) => 
                           X_Logic0_port, d(127) => X_Logic0_port, d(126) => 
                           X_Logic0_port, d(125) => X_Logic0_port, d(124) => 
                           X_Logic0_port, d(123) => X_Logic0_port, d(122) => 
                           X_Logic0_port, d(121) => X_Logic0_port, d(120) => 
                           X_Logic0_port, d(119) => X_Logic0_port, d(118) => 
                           X_Logic0_port, d(117) => X_Logic0_port, d(116) => 
                           X_Logic0_port, d(115) => X_Logic0_port, d(114) => 
                           X_Logic0_port, d(113) => X_Logic0_port, d(112) => 
                           X_Logic0_port, d(111) => X_Logic0_port, d(110) => 
                           X_Logic0_port, d(109) => X_Logic0_port, d(108) => 
                           X_Logic0_port, d(107) => X_Logic0_port, d(106) => 
                           X_Logic0_port, d(105) => X_Logic0_port, d(104) => 
                           X_Logic0_port, d(103) => X_Logic0_port, d(102) => 
                           X_Logic0_port, d(101) => X_Logic0_port, d(100) => 
                           X_Logic0_port, d(99) => X_Logic0_port, d(98) => 
                           muxes_in_4_150_port, d(97) => muxes_in_4_151_port, 
                           d(96) => muxes_in_4_152_port, d(95) => 
                           muxes_in_4_153_port, d(94) => muxes_in_4_154_port, 
                           d(93) => muxes_in_4_155_port, d(92) => 
                           muxes_in_4_156_port, d(91) => muxes_in_4_157_port, 
                           d(90) => muxes_in_4_158_port, d(89) => 
                           muxes_in_4_159_port, d(88) => muxes_in_4_160_port, 
                           d(87) => muxes_in_4_161_port, d(86) => 
                           muxes_in_4_162_port, d(85) => muxes_in_4_163_port, 
                           d(84) => muxes_in_4_164_port, d(83) => 
                           muxes_in_4_165_port, d(82) => muxes_in_4_166_port, 
                           d(81) => muxes_in_4_167_port, d(80) => 
                           muxes_in_4_168_port, d(79) => muxes_in_4_169_port, 
                           d(78) => muxes_in_4_170_port, d(77) => 
                           muxes_in_4_171_port, d(76) => muxes_in_4_172_port, 
                           d(75) => X_Logic0_port, d(74) => X_Logic0_port, 
                           d(73) => muxes_in_4_175_port, d(72) => 
                           muxes_in_4_176_port, d(71) => muxes_in_4_177_port, 
                           d(70) => muxes_in_4_178_port, d(69) => 
                           muxes_in_4_179_port, d(68) => muxes_in_4_180_port, 
                           d(67) => muxes_in_4_181_port, d(66) => 
                           muxes_in_4_182_port, d(65) => muxes_in_4_183_port, 
                           d(64) => muxes_in_4_184_port, d(63) => 
                           muxes_in_4_185_port, d(62) => muxes_in_4_186_port, 
                           d(61) => muxes_in_4_187_port, d(60) => 
                           muxes_in_4_188_port, d(59) => muxes_in_4_189_port, 
                           d(58) => muxes_in_4_190_port, d(57) => 
                           muxes_in_4_191_port, d(56) => muxes_in_4_192_port, 
                           d(55) => muxes_in_4_193_port, d(54) => 
                           muxes_in_4_194_port, d(53) => muxes_in_4_195_port, 
                           d(52) => muxes_in_4_196_port, d(51) => 
                           muxes_in_4_197_port, d(50) => X_Logic0_port, d(49) 
                           => X_Logic0_port, d(48) => X_Logic0_port, d(47) => 
                           X_Logic0_port, d(46) => X_Logic0_port, d(45) => 
                           X_Logic0_port, d(44) => X_Logic0_port, d(43) => 
                           X_Logic0_port, d(42) => X_Logic0_port, d(41) => 
                           X_Logic0_port, d(40) => X_Logic0_port, d(39) => 
                           X_Logic0_port, d(38) => X_Logic0_port, d(37) => 
                           X_Logic0_port, d(36) => X_Logic0_port, d(35) => 
                           X_Logic0_port, d(34) => X_Logic0_port, d(33) => 
                           X_Logic0_port, d(32) => X_Logic0_port, d(31) => 
                           X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           X_Logic0_port, d(20) => X_Logic0_port, d(19) => 
                           X_Logic0_port, d(18) => X_Logic0_port, d(17) => 
                           X_Logic0_port, d(16) => X_Logic0_port, d(15) => 
                           X_Logic0_port, d(14) => X_Logic0_port, d(13) => 
                           X_Logic0_port, d(12) => X_Logic0_port, d(11) => 
                           X_Logic0_port, d(10) => X_Logic0_port, d(9) => 
                           X_Logic0_port, d(8) => X_Logic0_port, d(7) => 
                           X_Logic0_port, d(6) => X_Logic0_port, d(5) => 
                           X_Logic0_port, d(4) => X_Logic0_port, d(3) => 
                           X_Logic0_port, d(2) => X_Logic0_port, d(1) => 
                           X_Logic0_port, d(0) => X_Logic0_port, Q(248) => 
                           n_3712, Q(247) => n_3713, Q(246) => n_3714, Q(245) 
                           => n_3715, Q(244) => n_3716, Q(243) => n_3717, 
                           Q(242) => n_3718, Q(241) => n_3719, Q(240) => n_3720
                           , Q(239) => n_3721, Q(238) => n_3722, Q(237) => 
                           n_3723, Q(236) => n_3724, Q(235) => n_3725, Q(234) 
                           => n_3726, Q(233) => n_3727, Q(232) => n_3728, 
                           Q(231) => n_3729, Q(230) => n_3730, Q(229) => n_3731
                           , Q(228) => n_3732, Q(227) => n_3733, Q(226) => 
                           n_3734, Q(225) => n_3735, Q(224) => n_3736, Q(223) 
                           => muxes_in_5_27_port, Q(222) => muxes_in_5_28_port,
                           Q(221) => muxes_in_5_29_port, Q(220) => 
                           muxes_in_5_30_port, Q(219) => muxes_in_5_31_port, 
                           Q(218) => muxes_in_5_32_port, Q(217) => 
                           muxes_in_5_33_port, Q(216) => muxes_in_5_34_port, 
                           Q(215) => muxes_in_5_35_port, Q(214) => 
                           muxes_in_5_36_port, Q(213) => muxes_in_5_37_port, 
                           Q(212) => muxes_in_5_38_port, Q(211) => 
                           muxes_in_5_39_port, Q(210) => muxes_in_5_40_port, 
                           Q(209) => muxes_in_5_41_port, Q(208) => 
                           muxes_in_5_42_port, Q(207) => muxes_in_5_43_port, 
                           Q(206) => muxes_in_5_44_port, Q(205) => 
                           muxes_in_5_45_port, Q(204) => muxes_in_5_46_port, 
                           Q(203) => muxes_in_5_47_port, Q(202) => 
                           muxes_in_5_48_port, Q(201) => muxes_in_5_49_port, 
                           Q(200) => muxes_in_5_50_port, Q(199) => 
                           muxes_in_5_51_port, Q(198) => muxes_in_5_54_port, 
                           Q(197) => muxes_in_5_55_port, Q(196) => 
                           muxes_in_5_56_port, Q(195) => muxes_in_5_57_port, 
                           Q(194) => muxes_in_5_58_port, Q(193) => 
                           muxes_in_5_59_port, Q(192) => muxes_in_5_60_port, 
                           Q(191) => muxes_in_5_61_port, Q(190) => 
                           muxes_in_5_62_port, Q(189) => muxes_in_5_63_port, 
                           Q(188) => muxes_in_5_64_port, Q(187) => 
                           muxes_in_5_65_port, Q(186) => muxes_in_5_66_port, 
                           Q(185) => muxes_in_5_67_port, Q(184) => 
                           muxes_in_5_68_port, Q(183) => muxes_in_5_69_port, 
                           Q(182) => muxes_in_5_70_port, Q(181) => 
                           muxes_in_5_71_port, Q(180) => muxes_in_5_72_port, 
                           Q(179) => muxes_in_5_73_port, Q(178) => 
                           muxes_in_5_74_port, Q(177) => muxes_in_5_75_port, 
                           Q(176) => muxes_in_5_76_port, Q(175) => 
                           muxes_in_5_77_port, Q(174) => muxes_in_5_78_port, 
                           Q(173) => n_3737, Q(172) => n_3738, Q(171) => n_3739
                           , Q(170) => n_3740, Q(169) => n_3741, Q(168) => 
                           n_3742, Q(167) => n_3743, Q(166) => n_3744, Q(165) 
                           => n_3745, Q(164) => n_3746, Q(163) => n_3747, 
                           Q(162) => n_3748, Q(161) => n_3749, Q(160) => n_3750
                           , Q(159) => n_3751, Q(158) => n_3752, Q(157) => 
                           n_3753, Q(156) => n_3754, Q(155) => n_3755, Q(154) 
                           => n_3756, Q(153) => n_3757, Q(152) => n_3758, 
                           Q(151) => n_3759, Q(150) => n_3760, Q(149) => n_3761
                           , Q(148) => n_3762, Q(147) => n_3763, Q(146) => 
                           n_3764, Q(145) => n_3765, Q(144) => n_3766, Q(143) 
                           => n_3767, Q(142) => n_3768, Q(141) => n_3769, 
                           Q(140) => n_3770, Q(139) => n_3771, Q(138) => n_3772
                           , Q(137) => n_3773, Q(136) => n_3774, Q(135) => 
                           n_3775, Q(134) => n_3776, Q(133) => n_3777, Q(132) 
                           => n_3778, Q(131) => n_3779, Q(130) => n_3780, 
                           Q(129) => n_3781, Q(128) => n_3782, Q(127) => n_3783
                           , Q(126) => n_3784, Q(125) => n_3785, Q(124) => 
                           n_3786, Q(123) => n_3787, Q(122) => n_3788, Q(121) 
                           => n_3789, Q(120) => n_3790, Q(119) => n_3791, 
                           Q(118) => n_3792, Q(117) => n_3793, Q(116) => n_3794
                           , Q(115) => n_3795, Q(114) => n_3796, Q(113) => 
                           n_3797, Q(112) => n_3798, Q(111) => n_3799, Q(110) 
                           => n_3800, Q(109) => n_3801, Q(108) => n_3802, 
                           Q(107) => n_3803, Q(106) => n_3804, Q(105) => n_3805
                           , Q(104) => n_3806, Q(103) => n_3807, Q(102) => 
                           n_3808, Q(101) => n_3809, Q(100) => n_3810, Q(99) =>
                           n_3811, Q(98) => muxes_in_5_162_port, Q(97) => 
                           muxes_in_5_163_port, Q(96) => muxes_in_5_164_port, 
                           Q(95) => muxes_in_5_165_port, Q(94) => 
                           muxes_in_5_166_port, Q(93) => muxes_in_5_167_port, 
                           Q(92) => muxes_in_5_168_port, Q(91) => 
                           muxes_in_5_169_port, Q(90) => muxes_in_5_170_port, 
                           Q(89) => muxes_in_5_171_port, Q(88) => 
                           muxes_in_5_172_port, Q(87) => muxes_in_5_173_port, 
                           Q(86) => muxes_in_5_174_port, Q(85) => 
                           muxes_in_5_175_port, Q(84) => muxes_in_5_176_port, 
                           Q(83) => muxes_in_5_177_port, Q(82) => 
                           muxes_in_5_178_port, Q(81) => muxes_in_5_179_port, 
                           Q(80) => muxes_in_5_180_port, Q(79) => 
                           muxes_in_5_181_port, Q(78) => muxes_in_5_182_port, 
                           Q(77) => muxes_in_5_183_port, Q(76) => 
                           muxes_in_5_184_port, Q(75) => muxes_in_5_185_port, 
                           Q(74) => muxes_in_5_186_port, Q(73) => 
                           muxes_in_5_189_port, Q(72) => muxes_in_5_190_port, 
                           Q(71) => muxes_in_5_191_port, Q(70) => 
                           muxes_in_5_192_port, Q(69) => muxes_in_5_193_port, 
                           Q(68) => muxes_in_5_194_port, Q(67) => 
                           muxes_in_5_195_port, Q(66) => muxes_in_5_196_port, 
                           Q(65) => muxes_in_5_197_port, Q(64) => 
                           muxes_in_5_198_port, Q(63) => muxes_in_5_199_port, 
                           Q(62) => muxes_in_5_200_port, Q(61) => 
                           muxes_in_5_201_port, Q(60) => muxes_in_5_202_port, 
                           Q(59) => muxes_in_5_203_port, Q(58) => 
                           muxes_in_5_204_port, Q(57) => muxes_in_5_205_port, 
                           Q(56) => muxes_in_5_206_port, Q(55) => 
                           muxes_in_5_207_port, Q(54) => muxes_in_5_208_port, 
                           Q(53) => muxes_in_5_209_port, Q(52) => 
                           muxes_in_5_210_port, Q(51) => muxes_in_5_211_port, 
                           Q(50) => muxes_in_5_212_port, Q(49) => 
                           muxes_in_5_213_port, Q(48) => n_3812, Q(47) => 
                           n_3813, Q(46) => n_3814, Q(45) => n_3815, Q(44) => 
                           n_3816, Q(43) => n_3817, Q(42) => n_3818, Q(41) => 
                           n_3819, Q(40) => n_3820, Q(39) => n_3821, Q(38) => 
                           n_3822, Q(37) => n_3823, Q(36) => n_3824, Q(35) => 
                           n_3825, Q(34) => n_3826, Q(33) => n_3827, Q(32) => 
                           n_3828, Q(31) => n_3829, Q(30) => n_3830, Q(29) => 
                           n_3831, Q(28) => n_3832, Q(27) => n_3833, Q(26) => 
                           n_3834, Q(25) => n_3835, Q(24) => n_3836, Q(23) => 
                           n_3837, Q(22) => n_3838, Q(21) => n_3839, Q(20) => 
                           n_3840, Q(19) => n_3841, Q(18) => n_3842, Q(17) => 
                           n_3843, Q(16) => n_3844, Q(15) => n_3845, Q(14) => 
                           n_3846, Q(13) => n_3847, Q(12) => n_3848, Q(11) => 
                           n_3849, Q(10) => n_3850, Q(9) => n_3851, Q(8) => 
                           n_3852, Q(7) => n_3853, Q(6) => n_3854, Q(5) => 
                           n_3855, Q(4) => n_3856, Q(3) => n_3857, Q(2) => 
                           n_3858, Q(1) => n_3859, Q(0) => n_3860);
   MUXi_4 : MUX_zbit_nbit_N25_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           X_Logic0_port, inputs(22) => X_Logic0_port, 
                           inputs(23) => X_Logic0_port, inputs(24) => 
                           X_Logic0_port, inputs(25) => muxes_in_4_25_port, 
                           inputs(26) => muxes_in_4_26_port, inputs(27) => 
                           muxes_in_4_27_port, inputs(28) => muxes_in_4_28_port
                           , inputs(29) => muxes_in_4_29_port, inputs(30) => 
                           muxes_in_4_30_port, inputs(31) => muxes_in_4_31_port
                           , inputs(32) => muxes_in_4_32_port, inputs(33) => 
                           muxes_in_4_33_port, inputs(34) => muxes_in_4_34_port
                           , inputs(35) => muxes_in_4_35_port, inputs(36) => 
                           muxes_in_4_36_port, inputs(37) => muxes_in_4_37_port
                           , inputs(38) => muxes_in_4_38_port, inputs(39) => 
                           muxes_in_4_39_port, inputs(40) => muxes_in_4_40_port
                           , inputs(41) => muxes_in_4_41_port, inputs(42) => 
                           muxes_in_4_42_port, inputs(43) => muxes_in_4_43_port
                           , inputs(44) => muxes_in_4_44_port, inputs(45) => 
                           muxes_in_4_45_port, inputs(46) => muxes_in_4_46_port
                           , inputs(47) => muxes_in_4_47_port, inputs(48) => 
                           X_Logic0_port, inputs(49) => X_Logic0_port, 
                           inputs(50) => muxes_in_4_50_port, inputs(51) => 
                           muxes_in_4_51_port, inputs(52) => muxes_in_4_52_port
                           , inputs(53) => muxes_in_4_53_port, inputs(54) => 
                           muxes_in_4_54_port, inputs(55) => muxes_in_4_55_port
                           , inputs(56) => muxes_in_4_56_port, inputs(57) => 
                           muxes_in_4_57_port, inputs(58) => muxes_in_4_58_port
                           , inputs(59) => muxes_in_4_59_port, inputs(60) => 
                           muxes_in_4_60_port, inputs(61) => muxes_in_4_61_port
                           , inputs(62) => muxes_in_4_62_port, inputs(63) => 
                           muxes_in_4_63_port, inputs(64) => muxes_in_4_64_port
                           , inputs(65) => muxes_in_4_65_port, inputs(66) => 
                           muxes_in_4_66_port, inputs(67) => muxes_in_4_67_port
                           , inputs(68) => muxes_in_4_68_port, inputs(69) => 
                           muxes_in_4_69_port, inputs(70) => muxes_in_4_70_port
                           , inputs(71) => muxes_in_4_71_port, inputs(72) => 
                           muxes_in_4_72_port, inputs(73) => X_Logic0_port, 
                           inputs(74) => X_Logic0_port, inputs(75) => 
                           X_Logic0_port, inputs(76) => X_Logic0_port, 
                           inputs(77) => X_Logic0_port, inputs(78) => 
                           X_Logic0_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           X_Logic0_port, inputs(127) => X_Logic0_port, 
                           inputs(128) => X_Logic0_port, inputs(129) => 
                           X_Logic0_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => X_Logic0_port, 
                           inputs(134) => X_Logic0_port, inputs(135) => 
                           X_Logic0_port, inputs(136) => X_Logic0_port, 
                           inputs(137) => X_Logic0_port, inputs(138) => 
                           X_Logic0_port, inputs(139) => X_Logic0_port, 
                           inputs(140) => X_Logic0_port, inputs(141) => 
                           X_Logic0_port, inputs(142) => X_Logic0_port, 
                           inputs(143) => X_Logic0_port, inputs(144) => 
                           X_Logic0_port, inputs(145) => X_Logic0_port, 
                           inputs(146) => X_Logic0_port, inputs(147) => 
                           X_Logic0_port, inputs(148) => X_Logic0_port, 
                           inputs(149) => X_Logic0_port, inputs(150) => 
                           muxes_in_4_150_port, inputs(151) => 
                           muxes_in_4_151_port, inputs(152) => 
                           muxes_in_4_152_port, inputs(153) => 
                           muxes_in_4_153_port, inputs(154) => 
                           muxes_in_4_154_port, inputs(155) => 
                           muxes_in_4_155_port, inputs(156) => 
                           muxes_in_4_156_port, inputs(157) => 
                           muxes_in_4_157_port, inputs(158) => 
                           muxes_in_4_158_port, inputs(159) => 
                           muxes_in_4_159_port, inputs(160) => 
                           muxes_in_4_160_port, inputs(161) => 
                           muxes_in_4_161_port, inputs(162) => 
                           muxes_in_4_162_port, inputs(163) => 
                           muxes_in_4_163_port, inputs(164) => 
                           muxes_in_4_164_port, inputs(165) => 
                           muxes_in_4_165_port, inputs(166) => 
                           muxes_in_4_166_port, inputs(167) => 
                           muxes_in_4_167_port, inputs(168) => 
                           muxes_in_4_168_port, inputs(169) => 
                           muxes_in_4_169_port, inputs(170) => 
                           muxes_in_4_170_port, inputs(171) => 
                           muxes_in_4_171_port, inputs(172) => 
                           muxes_in_4_172_port, inputs(173) => X_Logic0_port, 
                           inputs(174) => X_Logic0_port, inputs(175) => 
                           muxes_in_4_175_port, inputs(176) => 
                           muxes_in_4_176_port, inputs(177) => 
                           muxes_in_4_177_port, inputs(178) => 
                           muxes_in_4_178_port, inputs(179) => 
                           muxes_in_4_179_port, inputs(180) => 
                           muxes_in_4_180_port, inputs(181) => 
                           muxes_in_4_181_port, inputs(182) => 
                           muxes_in_4_182_port, inputs(183) => 
                           muxes_in_4_183_port, inputs(184) => 
                           muxes_in_4_184_port, inputs(185) => 
                           muxes_in_4_185_port, inputs(186) => 
                           muxes_in_4_186_port, inputs(187) => 
                           muxes_in_4_187_port, inputs(188) => 
                           muxes_in_4_188_port, inputs(189) => 
                           muxes_in_4_189_port, inputs(190) => 
                           muxes_in_4_190_port, inputs(191) => 
                           muxes_in_4_191_port, inputs(192) => 
                           muxes_in_4_192_port, inputs(193) => 
                           muxes_in_4_193_port, inputs(194) => 
                           muxes_in_4_194_port, inputs(195) => 
                           muxes_in_4_195_port, inputs(196) => 
                           muxes_in_4_196_port, inputs(197) => 
                           muxes_in_4_197_port, inputs(198) => X_Logic0_port, 
                           inputs(199) => X_Logic0_port, SEL(2) => 
                           encoder_out_4_2_port, SEL(1) => encoder_out_4_1_port
                           , SEL(0) => encoder_out_4_0_port, Y(24) => 
                           mux_out_4_24_port, Y(23) => mux_out_4_23_port, Y(22)
                           => mux_out_4_22_port, Y(21) => mux_out_4_21_port, 
                           Y(20) => mux_out_4_20_port, Y(19) => 
                           mux_out_4_19_port, Y(18) => mux_out_4_18_port, Y(17)
                           => mux_out_4_17_port, Y(16) => mux_out_4_16_port, 
                           Y(15) => mux_out_4_15_port, Y(14) => 
                           mux_out_4_14_port, Y(13) => mux_out_4_13_port, Y(12)
                           => mux_out_4_12_port, Y(11) => mux_out_4_11_port, 
                           Y(10) => mux_out_4_10_port, Y(9) => mux_out_4_9_port
                           , Y(8) => mux_out_4_8_port, Y(7) => mux_out_4_7_port
                           , Y(6) => mux_out_4_6_port, Y(5) => mux_out_4_5_port
                           , Y(4) => mux_out_4_4_port, Y(3) => mux_out_4_3_port
                           , Y(2) => mux_out_4_2_port, Y(1) => mux_out_4_1_port
                           , Y(0) => mux_out_4_0_port);
   ADDi_4 : adder_NBIT25 port map( a(24) => mux_out_4_24_port, a(23) => 
                           mux_out_4_23_port, a(22) => mux_out_4_22_port, a(21)
                           => mux_out_4_21_port, a(20) => mux_out_4_20_port, 
                           a(19) => mux_out_4_19_port, a(18) => 
                           mux_out_4_18_port, a(17) => mux_out_4_17_port, a(16)
                           => mux_out_4_16_port, a(15) => mux_out_4_15_port, 
                           a(14) => mux_out_4_14_port, a(13) => 
                           mux_out_4_13_port, a(12) => mux_out_4_12_port, a(11)
                           => mux_out_4_11_port, a(10) => mux_out_4_10_port, 
                           a(9) => mux_out_4_9_port, a(8) => mux_out_4_8_port, 
                           a(7) => mux_out_4_7_port, a(6) => mux_out_4_6_port, 
                           a(5) => mux_out_4_5_port, a(4) => mux_out_4_4_port, 
                           a(3) => mux_out_4_3_port, a(2) => mux_out_4_2_port, 
                           a(1) => mux_out_4_1_port, a(0) => mux_out_4_0_port, 
                           b(24) => sum_B_in_4_24_port, b(23) => 
                           sum_B_in_4_24_port, b(22) => sum_B_in_4_24_port, 
                           b(21) => sum_B_in_4_21_port, b(20) => 
                           sum_B_in_4_20_port, b(19) => sum_B_in_4_19_port, 
                           b(18) => sum_B_in_4_18_port, b(17) => 
                           sum_B_in_4_17_port, b(16) => sum_B_in_4_16_port, 
                           b(15) => sum_B_in_4_15_port, b(14) => 
                           sum_B_in_4_14_port, b(13) => sum_B_in_4_13_port, 
                           b(12) => sum_B_in_4_12_port, b(11) => 
                           sum_B_in_4_11_port, b(10) => sum_B_in_4_10_port, 
                           b(9) => sum_B_in_4_9_port, b(8) => sum_B_in_4_8_port
                           , b(7) => sum_B_in_4_7_port, b(6) => 
                           sum_B_in_4_6_port, b(5) => sum_B_in_4_5_port, b(4) 
                           => sum_B_in_4_4_port, b(3) => sum_B_in_4_3_port, 
                           b(2) => sum_B_in_4_2_port, b(1) => sum_B_in_4_1_port
                           , b(0) => sum_B_in_4_0_port, cin => X_Logic0_port, 
                           s(25) => sum_out_4_25_port, s(24) => 
                           sum_out_4_24_port, s(23) => sum_out_4_23_port, s(22)
                           => sum_out_4_22_port, s(21) => sum_out_4_21_port, 
                           s(20) => sum_out_4_20_port, s(19) => 
                           sum_out_4_19_port, s(18) => sum_out_4_18_port, s(17)
                           => sum_out_4_17_port, s(16) => sum_out_4_16_port, 
                           s(15) => sum_out_4_15_port, s(14) => 
                           sum_out_4_14_port, s(13) => sum_out_4_13_port, s(12)
                           => sum_out_4_12_port, s(11) => sum_out_4_11_port, 
                           s(10) => sum_out_4_10_port, s(9) => sum_out_4_9_port
                           , s(8) => sum_out_4_8_port, s(7) => sum_out_4_7_port
                           , s(6) => sum_out_4_6_port, s(5) => sum_out_4_5_port
                           , s(4) => sum_out_4_4_port, s(3) => sum_out_4_3_port
                           , s(2) => sum_out_4_2_port, s(1) => sum_out_4_1_port
                           , s(0) => sum_out_4_0_port);
   pip_del_reg_addi_4 : reg_nbit_n32_3 port map( clk => n12, reset => n6, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           sum_out_4_25_port, d(24) => sum_out_4_24_port, d(23)
                           => sum_out_4_23_port, d(22) => sum_out_4_22_port, 
                           d(21) => sum_out_4_21_port, d(20) => 
                           sum_out_4_20_port, d(19) => sum_out_4_19_port, d(18)
                           => sum_out_4_18_port, d(17) => sum_out_4_17_port, 
                           d(16) => sum_out_4_16_port, d(15) => 
                           sum_out_4_15_port, d(14) => sum_out_4_14_port, d(13)
                           => sum_out_4_13_port, d(12) => sum_out_4_12_port, 
                           d(11) => sum_out_4_11_port, d(10) => 
                           sum_out_4_10_port, d(9) => sum_out_4_9_port, d(8) =>
                           sum_out_4_8_port, d(7) => sum_out_4_7_port, d(6) => 
                           sum_out_4_6_port, d(5) => sum_out_4_5_port, d(4) => 
                           sum_out_4_4_port, d(3) => sum_out_4_3_port, d(2) => 
                           sum_out_4_2_port, d(1) => sum_out_4_1_port, d(0) => 
                           sum_out_4_0_port, Q(31) => n_3861, Q(30) => n_3862, 
                           Q(29) => n_3863, Q(28) => n_3864, Q(27) => n_3865, 
                           Q(26) => n_3866, Q(25) => n_3867, Q(24) => 
                           sum_B_in_5_26_port, Q(23) => sum_B_in_5_23_port, 
                           Q(22) => sum_B_in_5_22_port, Q(21) => 
                           sum_B_in_5_21_port, Q(20) => sum_B_in_5_20_port, 
                           Q(19) => sum_B_in_5_19_port, Q(18) => 
                           sum_B_in_5_18_port, Q(17) => sum_B_in_5_17_port, 
                           Q(16) => sum_B_in_5_16_port, Q(15) => 
                           sum_B_in_5_15_port, Q(14) => sum_B_in_5_14_port, 
                           Q(13) => sum_B_in_5_13_port, Q(12) => 
                           sum_B_in_5_12_port, Q(11) => sum_B_in_5_11_port, 
                           Q(10) => sum_B_in_5_10_port, Q(9) => 
                           sum_B_in_5_9_port, Q(8) => sum_B_in_5_8_port, Q(7) 
                           => sum_B_in_5_7_port, Q(6) => sum_B_in_5_6_port, 
                           Q(5) => sum_B_in_5_5_port, Q(4) => sum_B_in_5_4_port
                           , Q(3) => sum_B_in_5_3_port, Q(2) => 
                           sum_B_in_5_2_port, Q(1) => sum_B_in_5_1_port, Q(0) 
                           => sum_B_in_5_0_port);
   ENCi_5 : encoder_3 port map( y(2) => multiplicand_pip_5_11_port, y(1) => 
                           multiplicand_pip_5_10_port, y(0) => 
                           multiplicand_pip_5_9_port, sel(2) => 
                           encoder_out_5_2_port, sel(1) => encoder_out_5_1_port
                           , sel(0) => encoder_out_5_0_port);
   pip_del_reg_muxi_5 : reg_nbit_n249_3 port map( clk => n10, reset => n6, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => X_Logic0_port, 
                           d(226) => X_Logic0_port, d(225) => X_Logic0_port, 
                           d(224) => X_Logic0_port, d(223) => X_Logic0_port, 
                           d(222) => X_Logic0_port, d(221) => 
                           muxes_in_5_27_port, d(220) => muxes_in_5_28_port, 
                           d(219) => muxes_in_5_29_port, d(218) => 
                           muxes_in_5_30_port, d(217) => muxes_in_5_31_port, 
                           d(216) => muxes_in_5_32_port, d(215) => 
                           muxes_in_5_33_port, d(214) => muxes_in_5_34_port, 
                           d(213) => muxes_in_5_35_port, d(212) => 
                           muxes_in_5_36_port, d(211) => muxes_in_5_37_port, 
                           d(210) => muxes_in_5_38_port, d(209) => 
                           muxes_in_5_39_port, d(208) => muxes_in_5_40_port, 
                           d(207) => muxes_in_5_41_port, d(206) => 
                           muxes_in_5_42_port, d(205) => muxes_in_5_43_port, 
                           d(204) => muxes_in_5_44_port, d(203) => 
                           muxes_in_5_45_port, d(202) => muxes_in_5_46_port, 
                           d(201) => muxes_in_5_47_port, d(200) => 
                           muxes_in_5_48_port, d(199) => muxes_in_5_49_port, 
                           d(198) => muxes_in_5_50_port, d(197) => 
                           muxes_in_5_51_port, d(196) => X_Logic0_port, d(195) 
                           => X_Logic0_port, d(194) => muxes_in_5_54_port, 
                           d(193) => muxes_in_5_55_port, d(192) => 
                           muxes_in_5_56_port, d(191) => muxes_in_5_57_port, 
                           d(190) => muxes_in_5_58_port, d(189) => 
                           muxes_in_5_59_port, d(188) => muxes_in_5_60_port, 
                           d(187) => muxes_in_5_61_port, d(186) => 
                           muxes_in_5_62_port, d(185) => muxes_in_5_63_port, 
                           d(184) => muxes_in_5_64_port, d(183) => 
                           muxes_in_5_65_port, d(182) => muxes_in_5_66_port, 
                           d(181) => muxes_in_5_67_port, d(180) => 
                           muxes_in_5_68_port, d(179) => muxes_in_5_69_port, 
                           d(178) => muxes_in_5_70_port, d(177) => 
                           muxes_in_5_71_port, d(176) => muxes_in_5_72_port, 
                           d(175) => muxes_in_5_73_port, d(174) => 
                           muxes_in_5_74_port, d(173) => muxes_in_5_75_port, 
                           d(172) => muxes_in_5_76_port, d(171) => 
                           muxes_in_5_77_port, d(170) => muxes_in_5_78_port, 
                           d(169) => X_Logic0_port, d(168) => X_Logic0_port, 
                           d(167) => X_Logic0_port, d(166) => X_Logic0_port, 
                           d(165) => X_Logic0_port, d(164) => X_Logic0_port, 
                           d(163) => X_Logic0_port, d(162) => X_Logic0_port, 
                           d(161) => X_Logic0_port, d(160) => X_Logic0_port, 
                           d(159) => X_Logic0_port, d(158) => X_Logic0_port, 
                           d(157) => X_Logic0_port, d(156) => X_Logic0_port, 
                           d(155) => X_Logic0_port, d(154) => X_Logic0_port, 
                           d(153) => X_Logic0_port, d(152) => X_Logic0_port, 
                           d(151) => X_Logic0_port, d(150) => X_Logic0_port, 
                           d(149) => X_Logic0_port, d(148) => X_Logic0_port, 
                           d(147) => X_Logic0_port, d(146) => X_Logic0_port, 
                           d(145) => X_Logic0_port, d(144) => X_Logic0_port, 
                           d(143) => X_Logic0_port, d(142) => X_Logic0_port, 
                           d(141) => X_Logic0_port, d(140) => X_Logic0_port, 
                           d(139) => X_Logic0_port, d(138) => X_Logic0_port, 
                           d(137) => X_Logic0_port, d(136) => X_Logic0_port, 
                           d(135) => X_Logic0_port, d(134) => X_Logic0_port, 
                           d(133) => X_Logic0_port, d(132) => X_Logic0_port, 
                           d(131) => X_Logic0_port, d(130) => X_Logic0_port, 
                           d(129) => X_Logic0_port, d(128) => X_Logic0_port, 
                           d(127) => X_Logic0_port, d(126) => X_Logic0_port, 
                           d(125) => X_Logic0_port, d(124) => X_Logic0_port, 
                           d(123) => X_Logic0_port, d(122) => X_Logic0_port, 
                           d(121) => X_Logic0_port, d(120) => X_Logic0_port, 
                           d(119) => X_Logic0_port, d(118) => X_Logic0_port, 
                           d(117) => X_Logic0_port, d(116) => X_Logic0_port, 
                           d(115) => X_Logic0_port, d(114) => X_Logic0_port, 
                           d(113) => X_Logic0_port, d(112) => X_Logic0_port, 
                           d(111) => X_Logic0_port, d(110) => X_Logic0_port, 
                           d(109) => X_Logic0_port, d(108) => X_Logic0_port, 
                           d(107) => X_Logic0_port, d(106) => X_Logic0_port, 
                           d(105) => X_Logic0_port, d(104) => X_Logic0_port, 
                           d(103) => X_Logic0_port, d(102) => X_Logic0_port, 
                           d(101) => X_Logic0_port, d(100) => X_Logic0_port, 
                           d(99) => X_Logic0_port, d(98) => X_Logic0_port, 
                           d(97) => X_Logic0_port, d(96) => X_Logic0_port, 
                           d(95) => X_Logic0_port, d(94) => X_Logic0_port, 
                           d(93) => X_Logic0_port, d(92) => X_Logic0_port, 
                           d(91) => X_Logic0_port, d(90) => X_Logic0_port, 
                           d(89) => X_Logic0_port, d(88) => X_Logic0_port, 
                           d(87) => X_Logic0_port, d(86) => muxes_in_5_162_port
                           , d(85) => muxes_in_5_163_port, d(84) => 
                           muxes_in_5_164_port, d(83) => muxes_in_5_165_port, 
                           d(82) => muxes_in_5_166_port, d(81) => 
                           muxes_in_5_167_port, d(80) => muxes_in_5_168_port, 
                           d(79) => muxes_in_5_169_port, d(78) => 
                           muxes_in_5_170_port, d(77) => muxes_in_5_171_port, 
                           d(76) => muxes_in_5_172_port, d(75) => 
                           muxes_in_5_173_port, d(74) => muxes_in_5_174_port, 
                           d(73) => muxes_in_5_175_port, d(72) => 
                           muxes_in_5_176_port, d(71) => muxes_in_5_177_port, 
                           d(70) => muxes_in_5_178_port, d(69) => 
                           muxes_in_5_179_port, d(68) => muxes_in_5_180_port, 
                           d(67) => muxes_in_5_181_port, d(66) => 
                           muxes_in_5_182_port, d(65) => muxes_in_5_183_port, 
                           d(64) => muxes_in_5_184_port, d(63) => 
                           muxes_in_5_185_port, d(62) => muxes_in_5_186_port, 
                           d(61) => X_Logic0_port, d(60) => X_Logic0_port, 
                           d(59) => muxes_in_5_189_port, d(58) => 
                           muxes_in_5_190_port, d(57) => muxes_in_5_191_port, 
                           d(56) => muxes_in_5_192_port, d(55) => 
                           muxes_in_5_193_port, d(54) => muxes_in_5_194_port, 
                           d(53) => muxes_in_5_195_port, d(52) => 
                           muxes_in_5_196_port, d(51) => muxes_in_5_197_port, 
                           d(50) => muxes_in_5_198_port, d(49) => 
                           muxes_in_5_199_port, d(48) => muxes_in_5_200_port, 
                           d(47) => muxes_in_5_201_port, d(46) => 
                           muxes_in_5_202_port, d(45) => muxes_in_5_203_port, 
                           d(44) => muxes_in_5_204_port, d(43) => 
                           muxes_in_5_205_port, d(42) => muxes_in_5_206_port, 
                           d(41) => muxes_in_5_207_port, d(40) => 
                           muxes_in_5_208_port, d(39) => muxes_in_5_209_port, 
                           d(38) => muxes_in_5_210_port, d(37) => 
                           muxes_in_5_211_port, d(36) => muxes_in_5_212_port, 
                           d(35) => muxes_in_5_213_port, d(34) => X_Logic0_port
                           , d(33) => X_Logic0_port, d(32) => X_Logic0_port, 
                           d(31) => X_Logic0_port, d(30) => X_Logic0_port, 
                           d(29) => X_Logic0_port, d(28) => X_Logic0_port, 
                           d(27) => X_Logic0_port, d(26) => X_Logic0_port, 
                           d(25) => X_Logic0_port, d(24) => X_Logic0_port, 
                           d(23) => X_Logic0_port, d(22) => X_Logic0_port, 
                           d(21) => X_Logic0_port, d(20) => X_Logic0_port, 
                           d(19) => X_Logic0_port, d(18) => X_Logic0_port, 
                           d(17) => X_Logic0_port, d(16) => X_Logic0_port, 
                           d(15) => X_Logic0_port, d(14) => X_Logic0_port, 
                           d(13) => X_Logic0_port, d(12) => X_Logic0_port, 
                           d(11) => X_Logic0_port, d(10) => X_Logic0_port, d(9)
                           => X_Logic0_port, d(8) => X_Logic0_port, d(7) => 
                           X_Logic0_port, d(6) => X_Logic0_port, d(5) => 
                           X_Logic0_port, d(4) => X_Logic0_port, d(3) => 
                           X_Logic0_port, d(2) => X_Logic0_port, d(1) => 
                           X_Logic0_port, d(0) => X_Logic0_port, Q(248) => 
                           n_3868, Q(247) => n_3869, Q(246) => n_3870, Q(245) 
                           => n_3871, Q(244) => n_3872, Q(243) => n_3873, 
                           Q(242) => n_3874, Q(241) => n_3875, Q(240) => n_3876
                           , Q(239) => n_3877, Q(238) => n_3878, Q(237) => 
                           n_3879, Q(236) => n_3880, Q(235) => n_3881, Q(234) 
                           => n_3882, Q(233) => n_3883, Q(232) => n_3884, 
                           Q(231) => n_3885, Q(230) => n_3886, Q(229) => n_3887
                           , Q(228) => n_3888, Q(227) => n_3889, Q(226) => 
                           n_3890, Q(225) => n_3891, Q(224) => n_3892, Q(223) 
                           => n_3893, Q(222) => n_3894, Q(221) => 
                           muxes_in_6_29_port, Q(220) => muxes_in_6_30_port, 
                           Q(219) => muxes_in_6_31_port, Q(218) => 
                           muxes_in_6_32_port, Q(217) => muxes_in_6_33_port, 
                           Q(216) => muxes_in_6_34_port, Q(215) => 
                           muxes_in_6_35_port, Q(214) => muxes_in_6_36_port, 
                           Q(213) => muxes_in_6_37_port, Q(212) => 
                           muxes_in_6_38_port, Q(211) => muxes_in_6_39_port, 
                           Q(210) => muxes_in_6_40_port, Q(209) => 
                           muxes_in_6_41_port, Q(208) => muxes_in_6_42_port, 
                           Q(207) => muxes_in_6_43_port, Q(206) => 
                           muxes_in_6_44_port, Q(205) => muxes_in_6_45_port, 
                           Q(204) => muxes_in_6_46_port, Q(203) => 
                           muxes_in_6_47_port, Q(202) => muxes_in_6_48_port, 
                           Q(201) => muxes_in_6_49_port, Q(200) => 
                           muxes_in_6_50_port, Q(199) => muxes_in_6_51_port, 
                           Q(198) => muxes_in_6_52_port, Q(197) => 
                           muxes_in_6_53_port, Q(196) => muxes_in_6_54_port, 
                           Q(195) => muxes_in_6_55_port, Q(194) => 
                           muxes_in_6_58_port, Q(193) => muxes_in_6_59_port, 
                           Q(192) => muxes_in_6_60_port, Q(191) => 
                           muxes_in_6_61_port, Q(190) => muxes_in_6_62_port, 
                           Q(189) => muxes_in_6_63_port, Q(188) => 
                           muxes_in_6_64_port, Q(187) => muxes_in_6_65_port, 
                           Q(186) => muxes_in_6_66_port, Q(185) => 
                           muxes_in_6_67_port, Q(184) => muxes_in_6_68_port, 
                           Q(183) => muxes_in_6_69_port, Q(182) => 
                           muxes_in_6_70_port, Q(181) => muxes_in_6_71_port, 
                           Q(180) => muxes_in_6_72_port, Q(179) => 
                           muxes_in_6_73_port, Q(178) => muxes_in_6_74_port, 
                           Q(177) => muxes_in_6_75_port, Q(176) => 
                           muxes_in_6_76_port, Q(175) => muxes_in_6_77_port, 
                           Q(174) => muxes_in_6_78_port, Q(173) => 
                           muxes_in_6_79_port, Q(172) => muxes_in_6_80_port, 
                           Q(171) => muxes_in_6_81_port, Q(170) => 
                           muxes_in_6_82_port, Q(169) => muxes_in_6_83_port, 
                           Q(168) => muxes_in_6_84_port, Q(167) => n_3895, 
                           Q(166) => n_3896, Q(165) => n_3897, Q(164) => n_3898
                           , Q(163) => n_3899, Q(162) => n_3900, Q(161) => 
                           n_3901, Q(160) => n_3902, Q(159) => n_3903, Q(158) 
                           => n_3904, Q(157) => n_3905, Q(156) => n_3906, 
                           Q(155) => n_3907, Q(154) => n_3908, Q(153) => n_3909
                           , Q(152) => n_3910, Q(151) => n_3911, Q(150) => 
                           n_3912, Q(149) => n_3913, Q(148) => n_3914, Q(147) 
                           => n_3915, Q(146) => n_3916, Q(145) => n_3917, 
                           Q(144) => n_3918, Q(143) => n_3919, Q(142) => n_3920
                           , Q(141) => n_3921, Q(140) => n_3922, Q(139) => 
                           n_3923, Q(138) => n_3924, Q(137) => n_3925, Q(136) 
                           => n_3926, Q(135) => n_3927, Q(134) => n_3928, 
                           Q(133) => n_3929, Q(132) => n_3930, Q(131) => n_3931
                           , Q(130) => n_3932, Q(129) => n_3933, Q(128) => 
                           n_3934, Q(127) => n_3935, Q(126) => n_3936, Q(125) 
                           => n_3937, Q(124) => n_3938, Q(123) => n_3939, 
                           Q(122) => n_3940, Q(121) => n_3941, Q(120) => n_3942
                           , Q(119) => n_3943, Q(118) => n_3944, Q(117) => 
                           n_3945, Q(116) => n_3946, Q(115) => n_3947, Q(114) 
                           => n_3948, Q(113) => n_3949, Q(112) => n_3950, 
                           Q(111) => n_3951, Q(110) => n_3952, Q(109) => n_3953
                           , Q(108) => n_3954, Q(107) => n_3955, Q(106) => 
                           n_3956, Q(105) => n_3957, Q(104) => n_3958, Q(103) 
                           => n_3959, Q(102) => n_3960, Q(101) => n_3961, 
                           Q(100) => n_3962, Q(99) => n_3963, Q(98) => n_3964, 
                           Q(97) => n_3965, Q(96) => n_3966, Q(95) => n_3967, 
                           Q(94) => n_3968, Q(93) => n_3969, Q(92) => n_3970, 
                           Q(91) => n_3971, Q(90) => n_3972, Q(89) => n_3973, 
                           Q(88) => n_3974, Q(87) => n_3975, Q(86) => 
                           muxes_in_6_174_port, Q(85) => muxes_in_6_175_port, 
                           Q(84) => muxes_in_6_176_port, Q(83) => 
                           muxes_in_6_177_port, Q(82) => muxes_in_6_178_port, 
                           Q(81) => muxes_in_6_179_port, Q(80) => 
                           muxes_in_6_180_port, Q(79) => muxes_in_6_181_port, 
                           Q(78) => muxes_in_6_182_port, Q(77) => 
                           muxes_in_6_183_port, Q(76) => muxes_in_6_184_port, 
                           Q(75) => muxes_in_6_185_port, Q(74) => 
                           muxes_in_6_186_port, Q(73) => muxes_in_6_187_port, 
                           Q(72) => muxes_in_6_188_port, Q(71) => 
                           muxes_in_6_189_port, Q(70) => muxes_in_6_190_port, 
                           Q(69) => muxes_in_6_191_port, Q(68) => 
                           muxes_in_6_192_port, Q(67) => muxes_in_6_193_port, 
                           Q(66) => muxes_in_6_194_port, Q(65) => 
                           muxes_in_6_195_port, Q(64) => muxes_in_6_196_port, 
                           Q(63) => muxes_in_6_197_port, Q(62) => 
                           muxes_in_6_198_port, Q(61) => muxes_in_6_199_port, 
                           Q(60) => muxes_in_6_200_port, Q(59) => 
                           muxes_in_6_203_port, Q(58) => muxes_in_6_204_port, 
                           Q(57) => muxes_in_6_205_port, Q(56) => 
                           muxes_in_6_206_port, Q(55) => muxes_in_6_207_port, 
                           Q(54) => muxes_in_6_208_port, Q(53) => 
                           muxes_in_6_209_port, Q(52) => muxes_in_6_210_port, 
                           Q(51) => muxes_in_6_211_port, Q(50) => 
                           muxes_in_6_212_port, Q(49) => muxes_in_6_213_port, 
                           Q(48) => muxes_in_6_214_port, Q(47) => 
                           muxes_in_6_215_port, Q(46) => muxes_in_6_216_port, 
                           Q(45) => muxes_in_6_217_port, Q(44) => 
                           muxes_in_6_218_port, Q(43) => muxes_in_6_219_port, 
                           Q(42) => muxes_in_6_220_port, Q(41) => 
                           muxes_in_6_221_port, Q(40) => muxes_in_6_222_port, 
                           Q(39) => muxes_in_6_223_port, Q(38) => 
                           muxes_in_6_224_port, Q(37) => muxes_in_6_225_port, 
                           Q(36) => muxes_in_6_226_port, Q(35) => 
                           muxes_in_6_227_port, Q(34) => muxes_in_6_228_port, 
                           Q(33) => muxes_in_6_229_port, Q(32) => n_3976, Q(31)
                           => n_3977, Q(30) => n_3978, Q(29) => n_3979, Q(28) 
                           => n_3980, Q(27) => n_3981, Q(26) => n_3982, Q(25) 
                           => n_3983, Q(24) => n_3984, Q(23) => n_3985, Q(22) 
                           => n_3986, Q(21) => n_3987, Q(20) => n_3988, Q(19) 
                           => n_3989, Q(18) => n_3990, Q(17) => n_3991, Q(16) 
                           => n_3992, Q(15) => n_3993, Q(14) => n_3994, Q(13) 
                           => n_3995, Q(12) => n_3996, Q(11) => n_3997, Q(10) 
                           => n_3998, Q(9) => n_3999, Q(8) => n_4000, Q(7) => 
                           n_4001, Q(6) => n_4002, Q(5) => n_4003, Q(4) => 
                           n_4004, Q(3) => n_4005, Q(2) => n_4006, Q(1) => 
                           n_4007, Q(0) => n_4008);
   MUXi_5 : MUX_zbit_nbit_N27_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           X_Logic0_port, inputs(22) => X_Logic0_port, 
                           inputs(23) => X_Logic0_port, inputs(24) => 
                           X_Logic0_port, inputs(25) => X_Logic0_port, 
                           inputs(26) => X_Logic0_port, inputs(27) => 
                           muxes_in_5_27_port, inputs(28) => muxes_in_5_28_port
                           , inputs(29) => muxes_in_5_29_port, inputs(30) => 
                           muxes_in_5_30_port, inputs(31) => muxes_in_5_31_port
                           , inputs(32) => muxes_in_5_32_port, inputs(33) => 
                           muxes_in_5_33_port, inputs(34) => muxes_in_5_34_port
                           , inputs(35) => muxes_in_5_35_port, inputs(36) => 
                           muxes_in_5_36_port, inputs(37) => muxes_in_5_37_port
                           , inputs(38) => muxes_in_5_38_port, inputs(39) => 
                           muxes_in_5_39_port, inputs(40) => muxes_in_5_40_port
                           , inputs(41) => muxes_in_5_41_port, inputs(42) => 
                           muxes_in_5_42_port, inputs(43) => muxes_in_5_43_port
                           , inputs(44) => muxes_in_5_44_port, inputs(45) => 
                           muxes_in_5_45_port, inputs(46) => muxes_in_5_46_port
                           , inputs(47) => muxes_in_5_47_port, inputs(48) => 
                           muxes_in_5_48_port, inputs(49) => muxes_in_5_49_port
                           , inputs(50) => muxes_in_5_50_port, inputs(51) => 
                           muxes_in_5_51_port, inputs(52) => X_Logic0_port, 
                           inputs(53) => X_Logic0_port, inputs(54) => 
                           muxes_in_5_54_port, inputs(55) => muxes_in_5_55_port
                           , inputs(56) => muxes_in_5_56_port, inputs(57) => 
                           muxes_in_5_57_port, inputs(58) => muxes_in_5_58_port
                           , inputs(59) => muxes_in_5_59_port, inputs(60) => 
                           muxes_in_5_60_port, inputs(61) => muxes_in_5_61_port
                           , inputs(62) => muxes_in_5_62_port, inputs(63) => 
                           muxes_in_5_63_port, inputs(64) => muxes_in_5_64_port
                           , inputs(65) => muxes_in_5_65_port, inputs(66) => 
                           muxes_in_5_66_port, inputs(67) => muxes_in_5_67_port
                           , inputs(68) => muxes_in_5_68_port, inputs(69) => 
                           muxes_in_5_69_port, inputs(70) => muxes_in_5_70_port
                           , inputs(71) => muxes_in_5_71_port, inputs(72) => 
                           muxes_in_5_72_port, inputs(73) => muxes_in_5_73_port
                           , inputs(74) => muxes_in_5_74_port, inputs(75) => 
                           muxes_in_5_75_port, inputs(76) => muxes_in_5_76_port
                           , inputs(77) => muxes_in_5_77_port, inputs(78) => 
                           muxes_in_5_78_port, inputs(79) => X_Logic0_port, 
                           inputs(80) => X_Logic0_port, inputs(81) => 
                           X_Logic0_port, inputs(82) => X_Logic0_port, 
                           inputs(83) => X_Logic0_port, inputs(84) => 
                           X_Logic0_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           X_Logic0_port, inputs(127) => X_Logic0_port, 
                           inputs(128) => X_Logic0_port, inputs(129) => 
                           X_Logic0_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => X_Logic0_port, 
                           inputs(134) => X_Logic0_port, inputs(135) => 
                           X_Logic0_port, inputs(136) => X_Logic0_port, 
                           inputs(137) => X_Logic0_port, inputs(138) => 
                           X_Logic0_port, inputs(139) => X_Logic0_port, 
                           inputs(140) => X_Logic0_port, inputs(141) => 
                           X_Logic0_port, inputs(142) => X_Logic0_port, 
                           inputs(143) => X_Logic0_port, inputs(144) => 
                           X_Logic0_port, inputs(145) => X_Logic0_port, 
                           inputs(146) => X_Logic0_port, inputs(147) => 
                           X_Logic0_port, inputs(148) => X_Logic0_port, 
                           inputs(149) => X_Logic0_port, inputs(150) => 
                           X_Logic0_port, inputs(151) => X_Logic0_port, 
                           inputs(152) => X_Logic0_port, inputs(153) => 
                           X_Logic0_port, inputs(154) => X_Logic0_port, 
                           inputs(155) => X_Logic0_port, inputs(156) => 
                           X_Logic0_port, inputs(157) => X_Logic0_port, 
                           inputs(158) => X_Logic0_port, inputs(159) => 
                           X_Logic0_port, inputs(160) => X_Logic0_port, 
                           inputs(161) => X_Logic0_port, inputs(162) => 
                           muxes_in_5_162_port, inputs(163) => 
                           muxes_in_5_163_port, inputs(164) => 
                           muxes_in_5_164_port, inputs(165) => 
                           muxes_in_5_165_port, inputs(166) => 
                           muxes_in_5_166_port, inputs(167) => 
                           muxes_in_5_167_port, inputs(168) => 
                           muxes_in_5_168_port, inputs(169) => 
                           muxes_in_5_169_port, inputs(170) => 
                           muxes_in_5_170_port, inputs(171) => 
                           muxes_in_5_171_port, inputs(172) => 
                           muxes_in_5_172_port, inputs(173) => 
                           muxes_in_5_173_port, inputs(174) => 
                           muxes_in_5_174_port, inputs(175) => 
                           muxes_in_5_175_port, inputs(176) => 
                           muxes_in_5_176_port, inputs(177) => 
                           muxes_in_5_177_port, inputs(178) => 
                           muxes_in_5_178_port, inputs(179) => 
                           muxes_in_5_179_port, inputs(180) => 
                           muxes_in_5_180_port, inputs(181) => 
                           muxes_in_5_181_port, inputs(182) => 
                           muxes_in_5_182_port, inputs(183) => 
                           muxes_in_5_183_port, inputs(184) => 
                           muxes_in_5_184_port, inputs(185) => 
                           muxes_in_5_185_port, inputs(186) => 
                           muxes_in_5_186_port, inputs(187) => X_Logic0_port, 
                           inputs(188) => X_Logic0_port, inputs(189) => 
                           muxes_in_5_189_port, inputs(190) => 
                           muxes_in_5_190_port, inputs(191) => 
                           muxes_in_5_191_port, inputs(192) => 
                           muxes_in_5_192_port, inputs(193) => 
                           muxes_in_5_193_port, inputs(194) => 
                           muxes_in_5_194_port, inputs(195) => 
                           muxes_in_5_195_port, inputs(196) => 
                           muxes_in_5_196_port, inputs(197) => 
                           muxes_in_5_197_port, inputs(198) => 
                           muxes_in_5_198_port, inputs(199) => 
                           muxes_in_5_199_port, inputs(200) => 
                           muxes_in_5_200_port, inputs(201) => 
                           muxes_in_5_201_port, inputs(202) => 
                           muxes_in_5_202_port, inputs(203) => 
                           muxes_in_5_203_port, inputs(204) => 
                           muxes_in_5_204_port, inputs(205) => 
                           muxes_in_5_205_port, inputs(206) => 
                           muxes_in_5_206_port, inputs(207) => 
                           muxes_in_5_207_port, inputs(208) => 
                           muxes_in_5_208_port, inputs(209) => 
                           muxes_in_5_209_port, inputs(210) => 
                           muxes_in_5_210_port, inputs(211) => 
                           muxes_in_5_211_port, inputs(212) => 
                           muxes_in_5_212_port, inputs(213) => 
                           muxes_in_5_213_port, inputs(214) => X_Logic0_port, 
                           inputs(215) => X_Logic0_port, SEL(2) => 
                           encoder_out_5_2_port, SEL(1) => encoder_out_5_1_port
                           , SEL(0) => encoder_out_5_0_port, Y(26) => 
                           mux_out_5_26_port, Y(25) => mux_out_5_25_port, Y(24)
                           => mux_out_5_24_port, Y(23) => mux_out_5_23_port, 
                           Y(22) => mux_out_5_22_port, Y(21) => 
                           mux_out_5_21_port, Y(20) => mux_out_5_20_port, Y(19)
                           => mux_out_5_19_port, Y(18) => mux_out_5_18_port, 
                           Y(17) => mux_out_5_17_port, Y(16) => 
                           mux_out_5_16_port, Y(15) => mux_out_5_15_port, Y(14)
                           => mux_out_5_14_port, Y(13) => mux_out_5_13_port, 
                           Y(12) => mux_out_5_12_port, Y(11) => 
                           mux_out_5_11_port, Y(10) => mux_out_5_10_port, Y(9) 
                           => mux_out_5_9_port, Y(8) => mux_out_5_8_port, Y(7) 
                           => mux_out_5_7_port, Y(6) => mux_out_5_6_port, Y(5) 
                           => mux_out_5_5_port, Y(4) => mux_out_5_4_port, Y(3) 
                           => mux_out_5_3_port, Y(2) => mux_out_5_2_port, Y(1) 
                           => mux_out_5_1_port, Y(0) => mux_out_5_0_port);
   ADDi_5 : adder_NBIT27 port map( a(26) => mux_out_5_26_port, a(25) => 
                           mux_out_5_25_port, a(24) => mux_out_5_24_port, a(23)
                           => mux_out_5_23_port, a(22) => mux_out_5_22_port, 
                           a(21) => mux_out_5_21_port, a(20) => 
                           mux_out_5_20_port, a(19) => mux_out_5_19_port, a(18)
                           => mux_out_5_18_port, a(17) => mux_out_5_17_port, 
                           a(16) => mux_out_5_16_port, a(15) => 
                           mux_out_5_15_port, a(14) => mux_out_5_14_port, a(13)
                           => mux_out_5_13_port, a(12) => mux_out_5_12_port, 
                           a(11) => mux_out_5_11_port, a(10) => 
                           mux_out_5_10_port, a(9) => mux_out_5_9_port, a(8) =>
                           mux_out_5_8_port, a(7) => mux_out_5_7_port, a(6) => 
                           mux_out_5_6_port, a(5) => mux_out_5_5_port, a(4) => 
                           mux_out_5_4_port, a(3) => mux_out_5_3_port, a(2) => 
                           mux_out_5_2_port, a(1) => mux_out_5_1_port, a(0) => 
                           mux_out_5_0_port, b(26) => sum_B_in_5_26_port, b(25)
                           => sum_B_in_5_26_port, b(24) => sum_B_in_5_26_port, 
                           b(23) => sum_B_in_5_23_port, b(22) => 
                           sum_B_in_5_22_port, b(21) => sum_B_in_5_21_port, 
                           b(20) => sum_B_in_5_20_port, b(19) => 
                           sum_B_in_5_19_port, b(18) => sum_B_in_5_18_port, 
                           b(17) => sum_B_in_5_17_port, b(16) => 
                           sum_B_in_5_16_port, b(15) => sum_B_in_5_15_port, 
                           b(14) => sum_B_in_5_14_port, b(13) => 
                           sum_B_in_5_13_port, b(12) => sum_B_in_5_12_port, 
                           b(11) => sum_B_in_5_11_port, b(10) => 
                           sum_B_in_5_10_port, b(9) => sum_B_in_5_9_port, b(8) 
                           => sum_B_in_5_8_port, b(7) => sum_B_in_5_7_port, 
                           b(6) => sum_B_in_5_6_port, b(5) => sum_B_in_5_5_port
                           , b(4) => sum_B_in_5_4_port, b(3) => 
                           sum_B_in_5_3_port, b(2) => sum_B_in_5_2_port, b(1) 
                           => sum_B_in_5_1_port, b(0) => sum_B_in_5_0_port, cin
                           => X_Logic0_port, s(27) => sum_out_5_27_port, s(26) 
                           => sum_out_5_26_port, s(25) => sum_out_5_25_port, 
                           s(24) => sum_out_5_24_port, s(23) => 
                           sum_out_5_23_port, s(22) => sum_out_5_22_port, s(21)
                           => sum_out_5_21_port, s(20) => sum_out_5_20_port, 
                           s(19) => sum_out_5_19_port, s(18) => 
                           sum_out_5_18_port, s(17) => sum_out_5_17_port, s(16)
                           => sum_out_5_16_port, s(15) => sum_out_5_15_port, 
                           s(14) => sum_out_5_14_port, s(13) => 
                           sum_out_5_13_port, s(12) => sum_out_5_12_port, s(11)
                           => sum_out_5_11_port, s(10) => sum_out_5_10_port, 
                           s(9) => sum_out_5_9_port, s(8) => sum_out_5_8_port, 
                           s(7) => sum_out_5_7_port, s(6) => sum_out_5_6_port, 
                           s(5) => sum_out_5_5_port, s(4) => sum_out_5_4_port, 
                           s(3) => sum_out_5_3_port, s(2) => sum_out_5_2_port, 
                           s(1) => sum_out_5_1_port, s(0) => sum_out_5_0_port);
   pip_del_reg_addi_5 : reg_nbit_n32_2 port map( clk => n12, reset => n5, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           sum_out_5_27_port, d(26) => sum_out_5_26_port, d(25)
                           => sum_out_5_25_port, d(24) => sum_out_5_24_port, 
                           d(23) => sum_out_5_23_port, d(22) => 
                           sum_out_5_22_port, d(21) => sum_out_5_21_port, d(20)
                           => sum_out_5_20_port, d(19) => sum_out_5_19_port, 
                           d(18) => sum_out_5_18_port, d(17) => 
                           sum_out_5_17_port, d(16) => sum_out_5_16_port, d(15)
                           => sum_out_5_15_port, d(14) => sum_out_5_14_port, 
                           d(13) => sum_out_5_13_port, d(12) => 
                           sum_out_5_12_port, d(11) => sum_out_5_11_port, d(10)
                           => sum_out_5_10_port, d(9) => sum_out_5_9_port, d(8)
                           => sum_out_5_8_port, d(7) => sum_out_5_7_port, d(6) 
                           => sum_out_5_6_port, d(5) => sum_out_5_5_port, d(4) 
                           => sum_out_5_4_port, d(3) => sum_out_5_3_port, d(2) 
                           => sum_out_5_2_port, d(1) => sum_out_5_1_port, d(0) 
                           => sum_out_5_0_port, Q(31) => n_4009, Q(30) => 
                           n_4010, Q(29) => n_4011, Q(28) => n_4012, Q(27) => 
                           n_4013, Q(26) => sum_B_in_6_28_port, Q(25) => 
                           sum_B_in_6_25_port, Q(24) => sum_B_in_6_24_port, 
                           Q(23) => sum_B_in_6_23_port, Q(22) => 
                           sum_B_in_6_22_port, Q(21) => sum_B_in_6_21_port, 
                           Q(20) => sum_B_in_6_20_port, Q(19) => 
                           sum_B_in_6_19_port, Q(18) => sum_B_in_6_18_port, 
                           Q(17) => sum_B_in_6_17_port, Q(16) => 
                           sum_B_in_6_16_port, Q(15) => sum_B_in_6_15_port, 
                           Q(14) => sum_B_in_6_14_port, Q(13) => 
                           sum_B_in_6_13_port, Q(12) => sum_B_in_6_12_port, 
                           Q(11) => sum_B_in_6_11_port, Q(10) => 
                           sum_B_in_6_10_port, Q(9) => sum_B_in_6_9_port, Q(8) 
                           => sum_B_in_6_8_port, Q(7) => sum_B_in_6_7_port, 
                           Q(6) => sum_B_in_6_6_port, Q(5) => sum_B_in_6_5_port
                           , Q(4) => sum_B_in_6_4_port, Q(3) => 
                           sum_B_in_6_3_port, Q(2) => sum_B_in_6_2_port, Q(1) 
                           => sum_B_in_6_1_port, Q(0) => sum_B_in_6_0_port);
   ENCi_6 : encoder_2 port map( y(2) => multiplicand_pip_6_13_port, y(1) => 
                           multiplicand_pip_6_12_port, y(0) => 
                           multiplicand_pip_6_11_port, sel(2) => 
                           encoder_out_6_2_port, sel(1) => encoder_out_6_1_port
                           , sel(0) => encoder_out_6_0_port);
   pip_del_reg_muxi_6 : reg_nbit_n249_2 port map( clk => n9, reset => n6, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => X_Logic0_port, 
                           d(226) => X_Logic0_port, d(225) => X_Logic0_port, 
                           d(224) => X_Logic0_port, d(223) => X_Logic0_port, 
                           d(222) => X_Logic0_port, d(221) => X_Logic0_port, 
                           d(220) => X_Logic0_port, d(219) => 
                           muxes_in_6_29_port, d(218) => muxes_in_6_30_port, 
                           d(217) => muxes_in_6_31_port, d(216) => 
                           muxes_in_6_32_port, d(215) => muxes_in_6_33_port, 
                           d(214) => muxes_in_6_34_port, d(213) => 
                           muxes_in_6_35_port, d(212) => muxes_in_6_36_port, 
                           d(211) => muxes_in_6_37_port, d(210) => 
                           muxes_in_6_38_port, d(209) => muxes_in_6_39_port, 
                           d(208) => muxes_in_6_40_port, d(207) => 
                           muxes_in_6_41_port, d(206) => muxes_in_6_42_port, 
                           d(205) => muxes_in_6_43_port, d(204) => 
                           muxes_in_6_44_port, d(203) => muxes_in_6_45_port, 
                           d(202) => muxes_in_6_46_port, d(201) => 
                           muxes_in_6_47_port, d(200) => muxes_in_6_48_port, 
                           d(199) => muxes_in_6_49_port, d(198) => 
                           muxes_in_6_50_port, d(197) => muxes_in_6_51_port, 
                           d(196) => muxes_in_6_52_port, d(195) => 
                           muxes_in_6_53_port, d(194) => muxes_in_6_54_port, 
                           d(193) => muxes_in_6_55_port, d(192) => 
                           X_Logic0_port, d(191) => X_Logic0_port, d(190) => 
                           muxes_in_6_58_port, d(189) => muxes_in_6_59_port, 
                           d(188) => muxes_in_6_60_port, d(187) => 
                           muxes_in_6_61_port, d(186) => muxes_in_6_62_port, 
                           d(185) => muxes_in_6_63_port, d(184) => 
                           muxes_in_6_64_port, d(183) => muxes_in_6_65_port, 
                           d(182) => muxes_in_6_66_port, d(181) => 
                           muxes_in_6_67_port, d(180) => muxes_in_6_68_port, 
                           d(179) => muxes_in_6_69_port, d(178) => 
                           muxes_in_6_70_port, d(177) => muxes_in_6_71_port, 
                           d(176) => muxes_in_6_72_port, d(175) => 
                           muxes_in_6_73_port, d(174) => muxes_in_6_74_port, 
                           d(173) => muxes_in_6_75_port, d(172) => 
                           muxes_in_6_76_port, d(171) => muxes_in_6_77_port, 
                           d(170) => muxes_in_6_78_port, d(169) => 
                           muxes_in_6_79_port, d(168) => muxes_in_6_80_port, 
                           d(167) => muxes_in_6_81_port, d(166) => 
                           muxes_in_6_82_port, d(165) => muxes_in_6_83_port, 
                           d(164) => muxes_in_6_84_port, d(163) => 
                           X_Logic0_port, d(162) => X_Logic0_port, d(161) => 
                           X_Logic0_port, d(160) => X_Logic0_port, d(159) => 
                           X_Logic0_port, d(158) => X_Logic0_port, d(157) => 
                           X_Logic0_port, d(156) => X_Logic0_port, d(155) => 
                           X_Logic0_port, d(154) => X_Logic0_port, d(153) => 
                           X_Logic0_port, d(152) => X_Logic0_port, d(151) => 
                           X_Logic0_port, d(150) => X_Logic0_port, d(149) => 
                           X_Logic0_port, d(148) => X_Logic0_port, d(147) => 
                           X_Logic0_port, d(146) => X_Logic0_port, d(145) => 
                           X_Logic0_port, d(144) => X_Logic0_port, d(143) => 
                           X_Logic0_port, d(142) => X_Logic0_port, d(141) => 
                           X_Logic0_port, d(140) => X_Logic0_port, d(139) => 
                           X_Logic0_port, d(138) => X_Logic0_port, d(137) => 
                           X_Logic0_port, d(136) => X_Logic0_port, d(135) => 
                           X_Logic0_port, d(134) => X_Logic0_port, d(133) => 
                           X_Logic0_port, d(132) => X_Logic0_port, d(131) => 
                           X_Logic0_port, d(130) => X_Logic0_port, d(129) => 
                           X_Logic0_port, d(128) => X_Logic0_port, d(127) => 
                           X_Logic0_port, d(126) => X_Logic0_port, d(125) => 
                           X_Logic0_port, d(124) => X_Logic0_port, d(123) => 
                           X_Logic0_port, d(122) => X_Logic0_port, d(121) => 
                           X_Logic0_port, d(120) => X_Logic0_port, d(119) => 
                           X_Logic0_port, d(118) => X_Logic0_port, d(117) => 
                           X_Logic0_port, d(116) => X_Logic0_port, d(115) => 
                           X_Logic0_port, d(114) => X_Logic0_port, d(113) => 
                           X_Logic0_port, d(112) => X_Logic0_port, d(111) => 
                           X_Logic0_port, d(110) => X_Logic0_port, d(109) => 
                           X_Logic0_port, d(108) => X_Logic0_port, d(107) => 
                           X_Logic0_port, d(106) => X_Logic0_port, d(105) => 
                           X_Logic0_port, d(104) => X_Logic0_port, d(103) => 
                           X_Logic0_port, d(102) => X_Logic0_port, d(101) => 
                           X_Logic0_port, d(100) => X_Logic0_port, d(99) => 
                           X_Logic0_port, d(98) => X_Logic0_port, d(97) => 
                           X_Logic0_port, d(96) => X_Logic0_port, d(95) => 
                           X_Logic0_port, d(94) => X_Logic0_port, d(93) => 
                           X_Logic0_port, d(92) => X_Logic0_port, d(91) => 
                           X_Logic0_port, d(90) => X_Logic0_port, d(89) => 
                           X_Logic0_port, d(88) => X_Logic0_port, d(87) => 
                           X_Logic0_port, d(86) => X_Logic0_port, d(85) => 
                           X_Logic0_port, d(84) => X_Logic0_port, d(83) => 
                           X_Logic0_port, d(82) => X_Logic0_port, d(81) => 
                           X_Logic0_port, d(80) => X_Logic0_port, d(79) => 
                           X_Logic0_port, d(78) => X_Logic0_port, d(77) => 
                           X_Logic0_port, d(76) => X_Logic0_port, d(75) => 
                           X_Logic0_port, d(74) => muxes_in_6_174_port, d(73) 
                           => muxes_in_6_175_port, d(72) => muxes_in_6_176_port
                           , d(71) => muxes_in_6_177_port, d(70) => 
                           muxes_in_6_178_port, d(69) => muxes_in_6_179_port, 
                           d(68) => muxes_in_6_180_port, d(67) => 
                           muxes_in_6_181_port, d(66) => muxes_in_6_182_port, 
                           d(65) => muxes_in_6_183_port, d(64) => 
                           muxes_in_6_184_port, d(63) => muxes_in_6_185_port, 
                           d(62) => muxes_in_6_186_port, d(61) => 
                           muxes_in_6_187_port, d(60) => muxes_in_6_188_port, 
                           d(59) => muxes_in_6_189_port, d(58) => 
                           muxes_in_6_190_port, d(57) => muxes_in_6_191_port, 
                           d(56) => muxes_in_6_192_port, d(55) => 
                           muxes_in_6_193_port, d(54) => muxes_in_6_194_port, 
                           d(53) => muxes_in_6_195_port, d(52) => 
                           muxes_in_6_196_port, d(51) => muxes_in_6_197_port, 
                           d(50) => muxes_in_6_198_port, d(49) => 
                           muxes_in_6_199_port, d(48) => muxes_in_6_200_port, 
                           d(47) => X_Logic0_port, d(46) => X_Logic0_port, 
                           d(45) => muxes_in_6_203_port, d(44) => 
                           muxes_in_6_204_port, d(43) => muxes_in_6_205_port, 
                           d(42) => muxes_in_6_206_port, d(41) => 
                           muxes_in_6_207_port, d(40) => muxes_in_6_208_port, 
                           d(39) => muxes_in_6_209_port, d(38) => 
                           muxes_in_6_210_port, d(37) => muxes_in_6_211_port, 
                           d(36) => muxes_in_6_212_port, d(35) => 
                           muxes_in_6_213_port, d(34) => muxes_in_6_214_port, 
                           d(33) => muxes_in_6_215_port, d(32) => 
                           muxes_in_6_216_port, d(31) => muxes_in_6_217_port, 
                           d(30) => muxes_in_6_218_port, d(29) => 
                           muxes_in_6_219_port, d(28) => muxes_in_6_220_port, 
                           d(27) => muxes_in_6_221_port, d(26) => 
                           muxes_in_6_222_port, d(25) => muxes_in_6_223_port, 
                           d(24) => muxes_in_6_224_port, d(23) => 
                           muxes_in_6_225_port, d(22) => muxes_in_6_226_port, 
                           d(21) => muxes_in_6_227_port, d(20) => 
                           muxes_in_6_228_port, d(19) => muxes_in_6_229_port, 
                           d(18) => X_Logic0_port, d(17) => X_Logic0_port, 
                           d(16) => X_Logic0_port, d(15) => X_Logic0_port, 
                           d(14) => X_Logic0_port, d(13) => X_Logic0_port, 
                           d(12) => X_Logic0_port, d(11) => X_Logic0_port, 
                           d(10) => X_Logic0_port, d(9) => X_Logic0_port, d(8) 
                           => X_Logic0_port, d(7) => X_Logic0_port, d(6) => 
                           X_Logic0_port, d(5) => X_Logic0_port, d(4) => 
                           X_Logic0_port, d(3) => X_Logic0_port, d(2) => 
                           X_Logic0_port, d(1) => X_Logic0_port, d(0) => 
                           X_Logic0_port, Q(248) => n_4014, Q(247) => n_4015, 
                           Q(246) => n_4016, Q(245) => n_4017, Q(244) => n_4018
                           , Q(243) => n_4019, Q(242) => n_4020, Q(241) => 
                           n_4021, Q(240) => n_4022, Q(239) => n_4023, Q(238) 
                           => n_4024, Q(237) => n_4025, Q(236) => n_4026, 
                           Q(235) => n_4027, Q(234) => n_4028, Q(233) => n_4029
                           , Q(232) => n_4030, Q(231) => n_4031, Q(230) => 
                           n_4032, Q(229) => n_4033, Q(228) => n_4034, Q(227) 
                           => n_4035, Q(226) => n_4036, Q(225) => n_4037, 
                           Q(224) => n_4038, Q(223) => n_4039, Q(222) => n_4040
                           , Q(221) => n_4041, Q(220) => n_4042, Q(219) => 
                           muxes_in_7_31_port, Q(218) => muxes_in_7_32_port, 
                           Q(217) => muxes_in_7_33_port, Q(216) => 
                           muxes_in_7_34_port, Q(215) => muxes_in_7_35_port, 
                           Q(214) => muxes_in_7_36_port, Q(213) => 
                           muxes_in_7_37_port, Q(212) => muxes_in_7_38_port, 
                           Q(211) => muxes_in_7_39_port, Q(210) => 
                           muxes_in_7_40_port, Q(209) => muxes_in_7_41_port, 
                           Q(208) => muxes_in_7_42_port, Q(207) => 
                           muxes_in_7_43_port, Q(206) => muxes_in_7_44_port, 
                           Q(205) => muxes_in_7_45_port, Q(204) => 
                           muxes_in_7_46_port, Q(203) => muxes_in_7_47_port, 
                           Q(202) => muxes_in_7_48_port, Q(201) => 
                           muxes_in_7_49_port, Q(200) => muxes_in_7_50_port, 
                           Q(199) => muxes_in_7_51_port, Q(198) => 
                           muxes_in_7_52_port, Q(197) => muxes_in_7_53_port, 
                           Q(196) => muxes_in_7_54_port, Q(195) => 
                           muxes_in_7_55_port, Q(194) => muxes_in_7_56_port, 
                           Q(193) => muxes_in_7_57_port, Q(192) => 
                           muxes_in_7_58_port, Q(191) => muxes_in_7_59_port, 
                           Q(190) => muxes_in_7_62_port, Q(189) => 
                           muxes_in_7_63_port, Q(188) => muxes_in_7_64_port, 
                           Q(187) => muxes_in_7_65_port, Q(186) => 
                           muxes_in_7_66_port, Q(185) => muxes_in_7_67_port, 
                           Q(184) => muxes_in_7_68_port, Q(183) => 
                           muxes_in_7_69_port, Q(182) => muxes_in_7_70_port, 
                           Q(181) => muxes_in_7_71_port, Q(180) => 
                           muxes_in_7_72_port, Q(179) => muxes_in_7_73_port, 
                           Q(178) => muxes_in_7_74_port, Q(177) => 
                           muxes_in_7_75_port, Q(176) => muxes_in_7_76_port, 
                           Q(175) => muxes_in_7_77_port, Q(174) => 
                           muxes_in_7_78_port, Q(173) => muxes_in_7_79_port, 
                           Q(172) => muxes_in_7_80_port, Q(171) => 
                           muxes_in_7_81_port, Q(170) => muxes_in_7_82_port, 
                           Q(169) => muxes_in_7_83_port, Q(168) => 
                           muxes_in_7_84_port, Q(167) => muxes_in_7_85_port, 
                           Q(166) => muxes_in_7_86_port, Q(165) => 
                           muxes_in_7_87_port, Q(164) => muxes_in_7_88_port, 
                           Q(163) => muxes_in_7_89_port, Q(162) => 
                           muxes_in_7_90_port, Q(161) => n_4043, Q(160) => 
                           n_4044, Q(159) => n_4045, Q(158) => n_4046, Q(157) 
                           => n_4047, Q(156) => n_4048, Q(155) => n_4049, 
                           Q(154) => n_4050, Q(153) => n_4051, Q(152) => n_4052
                           , Q(151) => n_4053, Q(150) => n_4054, Q(149) => 
                           n_4055, Q(148) => n_4056, Q(147) => n_4057, Q(146) 
                           => n_4058, Q(145) => n_4059, Q(144) => n_4060, 
                           Q(143) => n_4061, Q(142) => n_4062, Q(141) => n_4063
                           , Q(140) => n_4064, Q(139) => n_4065, Q(138) => 
                           n_4066, Q(137) => n_4067, Q(136) => n_4068, Q(135) 
                           => n_4069, Q(134) => n_4070, Q(133) => n_4071, 
                           Q(132) => n_4072, Q(131) => n_4073, Q(130) => n_4074
                           , Q(129) => n_4075, Q(128) => n_4076, Q(127) => 
                           n_4077, Q(126) => n_4078, Q(125) => n_4079, Q(124) 
                           => n_4080, Q(123) => n_4081, Q(122) => n_4082, 
                           Q(121) => n_4083, Q(120) => n_4084, Q(119) => n_4085
                           , Q(118) => n_4086, Q(117) => n_4087, Q(116) => 
                           n_4088, Q(115) => n_4089, Q(114) => n_4090, Q(113) 
                           => n_4091, Q(112) => n_4092, Q(111) => n_4093, 
                           Q(110) => n_4094, Q(109) => n_4095, Q(108) => n_4096
                           , Q(107) => n_4097, Q(106) => n_4098, Q(105) => 
                           n_4099, Q(104) => n_4100, Q(103) => n_4101, Q(102) 
                           => n_4102, Q(101) => n_4103, Q(100) => n_4104, Q(99)
                           => n_4105, Q(98) => n_4106, Q(97) => n_4107, Q(96) 
                           => n_4108, Q(95) => n_4109, Q(94) => n_4110, Q(93) 
                           => n_4111, Q(92) => n_4112, Q(91) => n_4113, Q(90) 
                           => n_4114, Q(89) => n_4115, Q(88) => n_4116, Q(87) 
                           => n_4117, Q(86) => n_4118, Q(85) => n_4119, Q(84) 
                           => n_4120, Q(83) => n_4121, Q(82) => n_4122, Q(81) 
                           => n_4123, Q(80) => n_4124, Q(79) => n_4125, Q(78) 
                           => n_4126, Q(77) => n_4127, Q(76) => n_4128, Q(75) 
                           => n_4129, Q(74) => muxes_in_7_186_port, Q(73) => 
                           muxes_in_7_187_port, Q(72) => muxes_in_7_188_port, 
                           Q(71) => muxes_in_7_189_port, Q(70) => 
                           muxes_in_7_190_port, Q(69) => muxes_in_7_191_port, 
                           Q(68) => muxes_in_7_192_port, Q(67) => 
                           muxes_in_7_193_port, Q(66) => muxes_in_7_194_port, 
                           Q(65) => muxes_in_7_195_port, Q(64) => 
                           muxes_in_7_196_port, Q(63) => muxes_in_7_197_port, 
                           Q(62) => muxes_in_7_198_port, Q(61) => 
                           muxes_in_7_199_port, Q(60) => muxes_in_7_200_port, 
                           Q(59) => muxes_in_7_201_port, Q(58) => 
                           muxes_in_7_202_port, Q(57) => muxes_in_7_203_port, 
                           Q(56) => muxes_in_7_204_port, Q(55) => 
                           muxes_in_7_205_port, Q(54) => muxes_in_7_206_port, 
                           Q(53) => muxes_in_7_207_port, Q(52) => 
                           muxes_in_7_208_port, Q(51) => muxes_in_7_209_port, 
                           Q(50) => muxes_in_7_210_port, Q(49) => 
                           muxes_in_7_211_port, Q(48) => muxes_in_7_212_port, 
                           Q(47) => muxes_in_7_213_port, Q(46) => 
                           muxes_in_7_214_port, Q(45) => muxes_in_7_217_port, 
                           Q(44) => muxes_in_7_218_port, Q(43) => 
                           muxes_in_7_219_port, Q(42) => muxes_in_7_220_port, 
                           Q(41) => muxes_in_7_221_port, Q(40) => 
                           muxes_in_7_222_port, Q(39) => muxes_in_7_223_port, 
                           Q(38) => muxes_in_7_224_port, Q(37) => 
                           muxes_in_7_225_port, Q(36) => muxes_in_7_226_port, 
                           Q(35) => muxes_in_7_227_port, Q(34) => 
                           muxes_in_7_228_port, Q(33) => muxes_in_7_229_port, 
                           Q(32) => muxes_in_7_230_port, Q(31) => 
                           muxes_in_7_231_port, Q(30) => muxes_in_7_232_port, 
                           Q(29) => muxes_in_7_233_port, Q(28) => 
                           muxes_in_7_234_port, Q(27) => muxes_in_7_235_port, 
                           Q(26) => muxes_in_7_236_port, Q(25) => 
                           muxes_in_7_237_port, Q(24) => muxes_in_7_238_port, 
                           Q(23) => muxes_in_7_239_port, Q(22) => 
                           muxes_in_7_240_port, Q(21) => muxes_in_7_241_port, 
                           Q(20) => muxes_in_7_242_port, Q(19) => 
                           muxes_in_7_243_port, Q(18) => muxes_in_7_244_port, 
                           Q(17) => muxes_in_7_245_port, Q(16) => n_4130, Q(15)
                           => n_4131, Q(14) => n_4132, Q(13) => n_4133, Q(12) 
                           => n_4134, Q(11) => n_4135, Q(10) => n_4136, Q(9) =>
                           n_4137, Q(8) => n_4138, Q(7) => n_4139, Q(6) => 
                           n_4140, Q(5) => n_4141, Q(4) => n_4142, Q(3) => 
                           n_4143, Q(2) => n_4144, Q(1) => n_4145, Q(0) => 
                           n_4146);
   MUXi_6 : MUX_zbit_nbit_N29_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           X_Logic0_port, inputs(22) => X_Logic0_port, 
                           inputs(23) => X_Logic0_port, inputs(24) => 
                           X_Logic0_port, inputs(25) => X_Logic0_port, 
                           inputs(26) => X_Logic0_port, inputs(27) => 
                           X_Logic0_port, inputs(28) => X_Logic0_port, 
                           inputs(29) => muxes_in_6_29_port, inputs(30) => 
                           muxes_in_6_30_port, inputs(31) => muxes_in_6_31_port
                           , inputs(32) => muxes_in_6_32_port, inputs(33) => 
                           muxes_in_6_33_port, inputs(34) => muxes_in_6_34_port
                           , inputs(35) => muxes_in_6_35_port, inputs(36) => 
                           muxes_in_6_36_port, inputs(37) => muxes_in_6_37_port
                           , inputs(38) => muxes_in_6_38_port, inputs(39) => 
                           muxes_in_6_39_port, inputs(40) => muxes_in_6_40_port
                           , inputs(41) => muxes_in_6_41_port, inputs(42) => 
                           muxes_in_6_42_port, inputs(43) => muxes_in_6_43_port
                           , inputs(44) => muxes_in_6_44_port, inputs(45) => 
                           muxes_in_6_45_port, inputs(46) => muxes_in_6_46_port
                           , inputs(47) => muxes_in_6_47_port, inputs(48) => 
                           muxes_in_6_48_port, inputs(49) => muxes_in_6_49_port
                           , inputs(50) => muxes_in_6_50_port, inputs(51) => 
                           muxes_in_6_51_port, inputs(52) => muxes_in_6_52_port
                           , inputs(53) => muxes_in_6_53_port, inputs(54) => 
                           muxes_in_6_54_port, inputs(55) => muxes_in_6_55_port
                           , inputs(56) => X_Logic0_port, inputs(57) => 
                           X_Logic0_port, inputs(58) => muxes_in_6_58_port, 
                           inputs(59) => muxes_in_6_59_port, inputs(60) => 
                           muxes_in_6_60_port, inputs(61) => muxes_in_6_61_port
                           , inputs(62) => muxes_in_6_62_port, inputs(63) => 
                           muxes_in_6_63_port, inputs(64) => muxes_in_6_64_port
                           , inputs(65) => muxes_in_6_65_port, inputs(66) => 
                           muxes_in_6_66_port, inputs(67) => muxes_in_6_67_port
                           , inputs(68) => muxes_in_6_68_port, inputs(69) => 
                           muxes_in_6_69_port, inputs(70) => muxes_in_6_70_port
                           , inputs(71) => muxes_in_6_71_port, inputs(72) => 
                           muxes_in_6_72_port, inputs(73) => muxes_in_6_73_port
                           , inputs(74) => muxes_in_6_74_port, inputs(75) => 
                           muxes_in_6_75_port, inputs(76) => muxes_in_6_76_port
                           , inputs(77) => muxes_in_6_77_port, inputs(78) => 
                           muxes_in_6_78_port, inputs(79) => muxes_in_6_79_port
                           , inputs(80) => muxes_in_6_80_port, inputs(81) => 
                           muxes_in_6_81_port, inputs(82) => muxes_in_6_82_port
                           , inputs(83) => muxes_in_6_83_port, inputs(84) => 
                           muxes_in_6_84_port, inputs(85) => X_Logic0_port, 
                           inputs(86) => X_Logic0_port, inputs(87) => 
                           X_Logic0_port, inputs(88) => X_Logic0_port, 
                           inputs(89) => X_Logic0_port, inputs(90) => 
                           X_Logic0_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           X_Logic0_port, inputs(127) => X_Logic0_port, 
                           inputs(128) => X_Logic0_port, inputs(129) => 
                           X_Logic0_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => X_Logic0_port, 
                           inputs(134) => X_Logic0_port, inputs(135) => 
                           X_Logic0_port, inputs(136) => X_Logic0_port, 
                           inputs(137) => X_Logic0_port, inputs(138) => 
                           X_Logic0_port, inputs(139) => X_Logic0_port, 
                           inputs(140) => X_Logic0_port, inputs(141) => 
                           X_Logic0_port, inputs(142) => X_Logic0_port, 
                           inputs(143) => X_Logic0_port, inputs(144) => 
                           X_Logic0_port, inputs(145) => X_Logic0_port, 
                           inputs(146) => X_Logic0_port, inputs(147) => 
                           X_Logic0_port, inputs(148) => X_Logic0_port, 
                           inputs(149) => X_Logic0_port, inputs(150) => 
                           X_Logic0_port, inputs(151) => X_Logic0_port, 
                           inputs(152) => X_Logic0_port, inputs(153) => 
                           X_Logic0_port, inputs(154) => X_Logic0_port, 
                           inputs(155) => X_Logic0_port, inputs(156) => 
                           X_Logic0_port, inputs(157) => X_Logic0_port, 
                           inputs(158) => X_Logic0_port, inputs(159) => 
                           X_Logic0_port, inputs(160) => X_Logic0_port, 
                           inputs(161) => X_Logic0_port, inputs(162) => 
                           X_Logic0_port, inputs(163) => X_Logic0_port, 
                           inputs(164) => X_Logic0_port, inputs(165) => 
                           X_Logic0_port, inputs(166) => X_Logic0_port, 
                           inputs(167) => X_Logic0_port, inputs(168) => 
                           X_Logic0_port, inputs(169) => X_Logic0_port, 
                           inputs(170) => X_Logic0_port, inputs(171) => 
                           X_Logic0_port, inputs(172) => X_Logic0_port, 
                           inputs(173) => X_Logic0_port, inputs(174) => 
                           muxes_in_6_174_port, inputs(175) => 
                           muxes_in_6_175_port, inputs(176) => 
                           muxes_in_6_176_port, inputs(177) => 
                           muxes_in_6_177_port, inputs(178) => 
                           muxes_in_6_178_port, inputs(179) => 
                           muxes_in_6_179_port, inputs(180) => 
                           muxes_in_6_180_port, inputs(181) => 
                           muxes_in_6_181_port, inputs(182) => 
                           muxes_in_6_182_port, inputs(183) => 
                           muxes_in_6_183_port, inputs(184) => 
                           muxes_in_6_184_port, inputs(185) => 
                           muxes_in_6_185_port, inputs(186) => 
                           muxes_in_6_186_port, inputs(187) => 
                           muxes_in_6_187_port, inputs(188) => 
                           muxes_in_6_188_port, inputs(189) => 
                           muxes_in_6_189_port, inputs(190) => 
                           muxes_in_6_190_port, inputs(191) => 
                           muxes_in_6_191_port, inputs(192) => 
                           muxes_in_6_192_port, inputs(193) => 
                           muxes_in_6_193_port, inputs(194) => 
                           muxes_in_6_194_port, inputs(195) => 
                           muxes_in_6_195_port, inputs(196) => 
                           muxes_in_6_196_port, inputs(197) => 
                           muxes_in_6_197_port, inputs(198) => 
                           muxes_in_6_198_port, inputs(199) => 
                           muxes_in_6_199_port, inputs(200) => 
                           muxes_in_6_200_port, inputs(201) => X_Logic0_port, 
                           inputs(202) => X_Logic0_port, inputs(203) => 
                           muxes_in_6_203_port, inputs(204) => 
                           muxes_in_6_204_port, inputs(205) => 
                           muxes_in_6_205_port, inputs(206) => 
                           muxes_in_6_206_port, inputs(207) => 
                           muxes_in_6_207_port, inputs(208) => 
                           muxes_in_6_208_port, inputs(209) => 
                           muxes_in_6_209_port, inputs(210) => 
                           muxes_in_6_210_port, inputs(211) => 
                           muxes_in_6_211_port, inputs(212) => 
                           muxes_in_6_212_port, inputs(213) => 
                           muxes_in_6_213_port, inputs(214) => 
                           muxes_in_6_214_port, inputs(215) => 
                           muxes_in_6_215_port, inputs(216) => 
                           muxes_in_6_216_port, inputs(217) => 
                           muxes_in_6_217_port, inputs(218) => 
                           muxes_in_6_218_port, inputs(219) => 
                           muxes_in_6_219_port, inputs(220) => 
                           muxes_in_6_220_port, inputs(221) => 
                           muxes_in_6_221_port, inputs(222) => 
                           muxes_in_6_222_port, inputs(223) => 
                           muxes_in_6_223_port, inputs(224) => 
                           muxes_in_6_224_port, inputs(225) => 
                           muxes_in_6_225_port, inputs(226) => 
                           muxes_in_6_226_port, inputs(227) => 
                           muxes_in_6_227_port, inputs(228) => 
                           muxes_in_6_228_port, inputs(229) => 
                           muxes_in_6_229_port, inputs(230) => X_Logic0_port, 
                           inputs(231) => X_Logic0_port, SEL(2) => 
                           encoder_out_6_2_port, SEL(1) => encoder_out_6_1_port
                           , SEL(0) => encoder_out_6_0_port, Y(28) => 
                           mux_out_6_28_port, Y(27) => mux_out_6_27_port, Y(26)
                           => mux_out_6_26_port, Y(25) => mux_out_6_25_port, 
                           Y(24) => mux_out_6_24_port, Y(23) => 
                           mux_out_6_23_port, Y(22) => mux_out_6_22_port, Y(21)
                           => mux_out_6_21_port, Y(20) => mux_out_6_20_port, 
                           Y(19) => mux_out_6_19_port, Y(18) => 
                           mux_out_6_18_port, Y(17) => mux_out_6_17_port, Y(16)
                           => mux_out_6_16_port, Y(15) => mux_out_6_15_port, 
                           Y(14) => mux_out_6_14_port, Y(13) => 
                           mux_out_6_13_port, Y(12) => mux_out_6_12_port, Y(11)
                           => mux_out_6_11_port, Y(10) => mux_out_6_10_port, 
                           Y(9) => mux_out_6_9_port, Y(8) => mux_out_6_8_port, 
                           Y(7) => mux_out_6_7_port, Y(6) => mux_out_6_6_port, 
                           Y(5) => mux_out_6_5_port, Y(4) => mux_out_6_4_port, 
                           Y(3) => mux_out_6_3_port, Y(2) => mux_out_6_2_port, 
                           Y(1) => mux_out_6_1_port, Y(0) => mux_out_6_0_port);
   ADDi_6 : adder_NBIT29 port map( a(28) => mux_out_6_28_port, a(27) => 
                           mux_out_6_27_port, a(26) => mux_out_6_26_port, a(25)
                           => mux_out_6_25_port, a(24) => mux_out_6_24_port, 
                           a(23) => mux_out_6_23_port, a(22) => 
                           mux_out_6_22_port, a(21) => mux_out_6_21_port, a(20)
                           => mux_out_6_20_port, a(19) => mux_out_6_19_port, 
                           a(18) => mux_out_6_18_port, a(17) => 
                           mux_out_6_17_port, a(16) => mux_out_6_16_port, a(15)
                           => mux_out_6_15_port, a(14) => mux_out_6_14_port, 
                           a(13) => mux_out_6_13_port, a(12) => 
                           mux_out_6_12_port, a(11) => mux_out_6_11_port, a(10)
                           => mux_out_6_10_port, a(9) => mux_out_6_9_port, a(8)
                           => mux_out_6_8_port, a(7) => mux_out_6_7_port, a(6) 
                           => mux_out_6_6_port, a(5) => mux_out_6_5_port, a(4) 
                           => mux_out_6_4_port, a(3) => mux_out_6_3_port, a(2) 
                           => mux_out_6_2_port, a(1) => mux_out_6_1_port, a(0) 
                           => mux_out_6_0_port, b(28) => sum_B_in_6_28_port, 
                           b(27) => sum_B_in_6_28_port, b(26) => 
                           sum_B_in_6_28_port, b(25) => sum_B_in_6_25_port, 
                           b(24) => sum_B_in_6_24_port, b(23) => 
                           sum_B_in_6_23_port, b(22) => sum_B_in_6_22_port, 
                           b(21) => sum_B_in_6_21_port, b(20) => 
                           sum_B_in_6_20_port, b(19) => sum_B_in_6_19_port, 
                           b(18) => sum_B_in_6_18_port, b(17) => 
                           sum_B_in_6_17_port, b(16) => sum_B_in_6_16_port, 
                           b(15) => sum_B_in_6_15_port, b(14) => 
                           sum_B_in_6_14_port, b(13) => sum_B_in_6_13_port, 
                           b(12) => sum_B_in_6_12_port, b(11) => 
                           sum_B_in_6_11_port, b(10) => sum_B_in_6_10_port, 
                           b(9) => sum_B_in_6_9_port, b(8) => sum_B_in_6_8_port
                           , b(7) => sum_B_in_6_7_port, b(6) => 
                           sum_B_in_6_6_port, b(5) => sum_B_in_6_5_port, b(4) 
                           => sum_B_in_6_4_port, b(3) => sum_B_in_6_3_port, 
                           b(2) => sum_B_in_6_2_port, b(1) => sum_B_in_6_1_port
                           , b(0) => sum_B_in_6_0_port, cin => X_Logic0_port, 
                           s(29) => sum_out_6_29_port, s(28) => 
                           sum_out_6_28_port, s(27) => sum_out_6_27_port, s(26)
                           => sum_out_6_26_port, s(25) => sum_out_6_25_port, 
                           s(24) => sum_out_6_24_port, s(23) => 
                           sum_out_6_23_port, s(22) => sum_out_6_22_port, s(21)
                           => sum_out_6_21_port, s(20) => sum_out_6_20_port, 
                           s(19) => sum_out_6_19_port, s(18) => 
                           sum_out_6_18_port, s(17) => sum_out_6_17_port, s(16)
                           => sum_out_6_16_port, s(15) => sum_out_6_15_port, 
                           s(14) => sum_out_6_14_port, s(13) => 
                           sum_out_6_13_port, s(12) => sum_out_6_12_port, s(11)
                           => sum_out_6_11_port, s(10) => sum_out_6_10_port, 
                           s(9) => sum_out_6_9_port, s(8) => sum_out_6_8_port, 
                           s(7) => sum_out_6_7_port, s(6) => sum_out_6_6_port, 
                           s(5) => sum_out_6_5_port, s(4) => sum_out_6_4_port, 
                           s(3) => sum_out_6_3_port, s(2) => sum_out_6_2_port, 
                           s(1) => sum_out_6_1_port, s(0) => sum_out_6_0_port);
   pip_del_reg_addi_6 : reg_nbit_n32_1 port map( clk => n12, reset => n6, d(31)
                           => X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           sum_out_6_29_port, d(28) => sum_out_6_28_port, d(27)
                           => sum_out_6_27_port, d(26) => sum_out_6_26_port, 
                           d(25) => sum_out_6_25_port, d(24) => 
                           sum_out_6_24_port, d(23) => sum_out_6_23_port, d(22)
                           => sum_out_6_22_port, d(21) => sum_out_6_21_port, 
                           d(20) => sum_out_6_20_port, d(19) => 
                           sum_out_6_19_port, d(18) => sum_out_6_18_port, d(17)
                           => sum_out_6_17_port, d(16) => sum_out_6_16_port, 
                           d(15) => sum_out_6_15_port, d(14) => 
                           sum_out_6_14_port, d(13) => sum_out_6_13_port, d(12)
                           => sum_out_6_12_port, d(11) => sum_out_6_11_port, 
                           d(10) => sum_out_6_10_port, d(9) => sum_out_6_9_port
                           , d(8) => sum_out_6_8_port, d(7) => sum_out_6_7_port
                           , d(6) => sum_out_6_6_port, d(5) => sum_out_6_5_port
                           , d(4) => sum_out_6_4_port, d(3) => sum_out_6_3_port
                           , d(2) => sum_out_6_2_port, d(1) => sum_out_6_1_port
                           , d(0) => sum_out_6_0_port, Q(31) => n_4147, Q(30) 
                           => n_4148, Q(29) => n_4149, Q(28) => 
                           sum_B_in_7_30_port, Q(27) => sum_B_in_7_27_port, 
                           Q(26) => sum_B_in_7_26_port, Q(25) => 
                           sum_B_in_7_25_port, Q(24) => sum_B_in_7_24_port, 
                           Q(23) => sum_B_in_7_23_port, Q(22) => 
                           sum_B_in_7_22_port, Q(21) => sum_B_in_7_21_port, 
                           Q(20) => sum_B_in_7_20_port, Q(19) => 
                           sum_B_in_7_19_port, Q(18) => sum_B_in_7_18_port, 
                           Q(17) => sum_B_in_7_17_port, Q(16) => 
                           sum_B_in_7_16_port, Q(15) => sum_B_in_7_15_port, 
                           Q(14) => sum_B_in_7_14_port, Q(13) => 
                           sum_B_in_7_13_port, Q(12) => sum_B_in_7_12_port, 
                           Q(11) => sum_B_in_7_11_port, Q(10) => 
                           sum_B_in_7_10_port, Q(9) => sum_B_in_7_9_port, Q(8) 
                           => sum_B_in_7_8_port, Q(7) => sum_B_in_7_7_port, 
                           Q(6) => sum_B_in_7_6_port, Q(5) => sum_B_in_7_5_port
                           , Q(4) => sum_B_in_7_4_port, Q(3) => 
                           sum_B_in_7_3_port, Q(2) => sum_B_in_7_2_port, Q(1) 
                           => sum_B_in_7_1_port, Q(0) => sum_B_in_7_0_port);
   ENCi_7 : encoder_1 port map( y(2) => multiplicand_pip_7_15_port, y(1) => 
                           multiplicand_pip_7_14_port, y(0) => 
                           multiplicand_pip_7_13_port, sel(2) => 
                           encoder_out_7_2_port, sel(1) => encoder_out_7_1_port
                           , sel(0) => encoder_out_7_0_port);
   pip_del_reg_muxi_7 : reg_nbit_n249_1 port map( clk => n9, reset => n5, 
                           d(248) => X_Logic0_port, d(247) => X_Logic0_port, 
                           d(246) => X_Logic0_port, d(245) => X_Logic0_port, 
                           d(244) => X_Logic0_port, d(243) => X_Logic0_port, 
                           d(242) => X_Logic0_port, d(241) => X_Logic0_port, 
                           d(240) => X_Logic0_port, d(239) => X_Logic0_port, 
                           d(238) => X_Logic0_port, d(237) => X_Logic0_port, 
                           d(236) => X_Logic0_port, d(235) => X_Logic0_port, 
                           d(234) => X_Logic0_port, d(233) => X_Logic0_port, 
                           d(232) => X_Logic0_port, d(231) => X_Logic0_port, 
                           d(230) => X_Logic0_port, d(229) => X_Logic0_port, 
                           d(228) => X_Logic0_port, d(227) => X_Logic0_port, 
                           d(226) => X_Logic0_port, d(225) => X_Logic0_port, 
                           d(224) => X_Logic0_port, d(223) => X_Logic0_port, 
                           d(222) => X_Logic0_port, d(221) => X_Logic0_port, 
                           d(220) => X_Logic0_port, d(219) => X_Logic0_port, 
                           d(218) => X_Logic0_port, d(217) => 
                           muxes_in_7_31_port, d(216) => muxes_in_7_32_port, 
                           d(215) => muxes_in_7_33_port, d(214) => 
                           muxes_in_7_34_port, d(213) => muxes_in_7_35_port, 
                           d(212) => muxes_in_7_36_port, d(211) => 
                           muxes_in_7_37_port, d(210) => muxes_in_7_38_port, 
                           d(209) => muxes_in_7_39_port, d(208) => 
                           muxes_in_7_40_port, d(207) => muxes_in_7_41_port, 
                           d(206) => muxes_in_7_42_port, d(205) => 
                           muxes_in_7_43_port, d(204) => muxes_in_7_44_port, 
                           d(203) => muxes_in_7_45_port, d(202) => 
                           muxes_in_7_46_port, d(201) => muxes_in_7_47_port, 
                           d(200) => muxes_in_7_48_port, d(199) => 
                           muxes_in_7_49_port, d(198) => muxes_in_7_50_port, 
                           d(197) => muxes_in_7_51_port, d(196) => 
                           muxes_in_7_52_port, d(195) => muxes_in_7_53_port, 
                           d(194) => muxes_in_7_54_port, d(193) => 
                           muxes_in_7_55_port, d(192) => muxes_in_7_56_port, 
                           d(191) => muxes_in_7_57_port, d(190) => 
                           muxes_in_7_58_port, d(189) => muxes_in_7_59_port, 
                           d(188) => X_Logic0_port, d(187) => X_Logic0_port, 
                           d(186) => muxes_in_7_62_port, d(185) => 
                           muxes_in_7_63_port, d(184) => muxes_in_7_64_port, 
                           d(183) => muxes_in_7_65_port, d(182) => 
                           muxes_in_7_66_port, d(181) => muxes_in_7_67_port, 
                           d(180) => muxes_in_7_68_port, d(179) => 
                           muxes_in_7_69_port, d(178) => muxes_in_7_70_port, 
                           d(177) => muxes_in_7_71_port, d(176) => 
                           muxes_in_7_72_port, d(175) => muxes_in_7_73_port, 
                           d(174) => muxes_in_7_74_port, d(173) => 
                           muxes_in_7_75_port, d(172) => muxes_in_7_76_port, 
                           d(171) => muxes_in_7_77_port, d(170) => 
                           muxes_in_7_78_port, d(169) => muxes_in_7_79_port, 
                           d(168) => muxes_in_7_80_port, d(167) => 
                           muxes_in_7_81_port, d(166) => muxes_in_7_82_port, 
                           d(165) => muxes_in_7_83_port, d(164) => 
                           muxes_in_7_84_port, d(163) => muxes_in_7_85_port, 
                           d(162) => muxes_in_7_86_port, d(161) => 
                           muxes_in_7_87_port, d(160) => muxes_in_7_88_port, 
                           d(159) => muxes_in_7_89_port, d(158) => 
                           muxes_in_7_90_port, d(157) => X_Logic0_port, d(156) 
                           => X_Logic0_port, d(155) => X_Logic0_port, d(154) =>
                           X_Logic0_port, d(153) => X_Logic0_port, d(152) => 
                           X_Logic0_port, d(151) => X_Logic0_port, d(150) => 
                           X_Logic0_port, d(149) => X_Logic0_port, d(148) => 
                           X_Logic0_port, d(147) => X_Logic0_port, d(146) => 
                           X_Logic0_port, d(145) => X_Logic0_port, d(144) => 
                           X_Logic0_port, d(143) => X_Logic0_port, d(142) => 
                           X_Logic0_port, d(141) => X_Logic0_port, d(140) => 
                           X_Logic0_port, d(139) => X_Logic0_port, d(138) => 
                           X_Logic0_port, d(137) => X_Logic0_port, d(136) => 
                           X_Logic0_port, d(135) => X_Logic0_port, d(134) => 
                           X_Logic0_port, d(133) => X_Logic0_port, d(132) => 
                           X_Logic0_port, d(131) => X_Logic0_port, d(130) => 
                           X_Logic0_port, d(129) => X_Logic0_port, d(128) => 
                           X_Logic0_port, d(127) => X_Logic0_port, d(126) => 
                           X_Logic0_port, d(125) => X_Logic0_port, d(124) => 
                           X_Logic0_port, d(123) => X_Logic0_port, d(122) => 
                           X_Logic0_port, d(121) => X_Logic0_port, d(120) => 
                           X_Logic0_port, d(119) => X_Logic0_port, d(118) => 
                           X_Logic0_port, d(117) => X_Logic0_port, d(116) => 
                           X_Logic0_port, d(115) => X_Logic0_port, d(114) => 
                           X_Logic0_port, d(113) => X_Logic0_port, d(112) => 
                           X_Logic0_port, d(111) => X_Logic0_port, d(110) => 
                           X_Logic0_port, d(109) => X_Logic0_port, d(108) => 
                           X_Logic0_port, d(107) => X_Logic0_port, d(106) => 
                           X_Logic0_port, d(105) => X_Logic0_port, d(104) => 
                           X_Logic0_port, d(103) => X_Logic0_port, d(102) => 
                           X_Logic0_port, d(101) => X_Logic0_port, d(100) => 
                           X_Logic0_port, d(99) => X_Logic0_port, d(98) => 
                           X_Logic0_port, d(97) => X_Logic0_port, d(96) => 
                           X_Logic0_port, d(95) => X_Logic0_port, d(94) => 
                           X_Logic0_port, d(93) => X_Logic0_port, d(92) => 
                           X_Logic0_port, d(91) => X_Logic0_port, d(90) => 
                           X_Logic0_port, d(89) => X_Logic0_port, d(88) => 
                           X_Logic0_port, d(87) => X_Logic0_port, d(86) => 
                           X_Logic0_port, d(85) => X_Logic0_port, d(84) => 
                           X_Logic0_port, d(83) => X_Logic0_port, d(82) => 
                           X_Logic0_port, d(81) => X_Logic0_port, d(80) => 
                           X_Logic0_port, d(79) => X_Logic0_port, d(78) => 
                           X_Logic0_port, d(77) => X_Logic0_port, d(76) => 
                           X_Logic0_port, d(75) => X_Logic0_port, d(74) => 
                           X_Logic0_port, d(73) => X_Logic0_port, d(72) => 
                           X_Logic0_port, d(71) => X_Logic0_port, d(70) => 
                           X_Logic0_port, d(69) => X_Logic0_port, d(68) => 
                           X_Logic0_port, d(67) => X_Logic0_port, d(66) => 
                           X_Logic0_port, d(65) => X_Logic0_port, d(64) => 
                           X_Logic0_port, d(63) => X_Logic0_port, d(62) => 
                           muxes_in_7_186_port, d(61) => muxes_in_7_187_port, 
                           d(60) => muxes_in_7_188_port, d(59) => 
                           muxes_in_7_189_port, d(58) => muxes_in_7_190_port, 
                           d(57) => muxes_in_7_191_port, d(56) => 
                           muxes_in_7_192_port, d(55) => muxes_in_7_193_port, 
                           d(54) => muxes_in_7_194_port, d(53) => 
                           muxes_in_7_195_port, d(52) => muxes_in_7_196_port, 
                           d(51) => muxes_in_7_197_port, d(50) => 
                           muxes_in_7_198_port, d(49) => muxes_in_7_199_port, 
                           d(48) => muxes_in_7_200_port, d(47) => 
                           muxes_in_7_201_port, d(46) => muxes_in_7_202_port, 
                           d(45) => muxes_in_7_203_port, d(44) => 
                           muxes_in_7_204_port, d(43) => muxes_in_7_205_port, 
                           d(42) => muxes_in_7_206_port, d(41) => 
                           muxes_in_7_207_port, d(40) => muxes_in_7_208_port, 
                           d(39) => muxes_in_7_209_port, d(38) => 
                           muxes_in_7_210_port, d(37) => muxes_in_7_211_port, 
                           d(36) => muxes_in_7_212_port, d(35) => 
                           muxes_in_7_213_port, d(34) => muxes_in_7_214_port, 
                           d(33) => X_Logic0_port, d(32) => X_Logic0_port, 
                           d(31) => muxes_in_7_217_port, d(30) => 
                           muxes_in_7_218_port, d(29) => muxes_in_7_219_port, 
                           d(28) => muxes_in_7_220_port, d(27) => 
                           muxes_in_7_221_port, d(26) => muxes_in_7_222_port, 
                           d(25) => muxes_in_7_223_port, d(24) => 
                           muxes_in_7_224_port, d(23) => muxes_in_7_225_port, 
                           d(22) => muxes_in_7_226_port, d(21) => 
                           muxes_in_7_227_port, d(20) => muxes_in_7_228_port, 
                           d(19) => muxes_in_7_229_port, d(18) => 
                           muxes_in_7_230_port, d(17) => muxes_in_7_231_port, 
                           d(16) => muxes_in_7_232_port, d(15) => 
                           muxes_in_7_233_port, d(14) => muxes_in_7_234_port, 
                           d(13) => muxes_in_7_235_port, d(12) => 
                           muxes_in_7_236_port, d(11) => muxes_in_7_237_port, 
                           d(10) => muxes_in_7_238_port, d(9) => 
                           muxes_in_7_239_port, d(8) => muxes_in_7_240_port, 
                           d(7) => muxes_in_7_241_port, d(6) => 
                           muxes_in_7_242_port, d(5) => muxes_in_7_243_port, 
                           d(4) => muxes_in_7_244_port, d(3) => 
                           muxes_in_7_245_port, d(2) => X_Logic0_port, d(1) => 
                           X_Logic0_port, d(0) => X_Logic0_port, Q(248) => 
                           n_4150, Q(247) => n_4151, Q(246) => n_4152, Q(245) 
                           => n_4153, Q(244) => n_4154, Q(243) => n_4155, 
                           Q(242) => n_4156, Q(241) => n_4157, Q(240) => n_4158
                           , Q(239) => n_4159, Q(238) => n_4160, Q(237) => 
                           n_4161, Q(236) => n_4162, Q(235) => n_4163, Q(234) 
                           => n_4164, Q(233) => n_4165, Q(232) => n_4166, 
                           Q(231) => n_4167, Q(230) => n_4168, Q(229) => n_4169
                           , Q(228) => n_4170, Q(227) => n_4171, Q(226) => 
                           n_4172, Q(225) => n_4173, Q(224) => n_4174, Q(223) 
                           => n_4175, Q(222) => n_4176, Q(221) => n_4177, 
                           Q(220) => n_4178, Q(219) => n_4179, Q(218) => n_4180
                           , Q(217) => n_4181, Q(216) => n_4182, Q(215) => 
                           n_4183, Q(214) => n_4184, Q(213) => n_4185, Q(212) 
                           => n_4186, Q(211) => n_4187, Q(210) => n_4188, 
                           Q(209) => n_4189, Q(208) => n_4190, Q(207) => n_4191
                           , Q(206) => n_4192, Q(205) => n_4193, Q(204) => 
                           n_4194, Q(203) => n_4195, Q(202) => n_4196, Q(201) 
                           => n_4197, Q(200) => n_4198, Q(199) => n_4199, 
                           Q(198) => n_4200, Q(197) => n_4201, Q(196) => n_4202
                           , Q(195) => n_4203, Q(194) => n_4204, Q(193) => 
                           n_4205, Q(192) => n_4206, Q(191) => n_4207, Q(190) 
                           => n_4208, Q(189) => n_4209, Q(188) => n_4210, 
                           Q(187) => n_4211, Q(186) => n_4212, Q(185) => n_4213
                           , Q(184) => n_4214, Q(183) => n_4215, Q(182) => 
                           n_4216, Q(181) => n_4217, Q(180) => n_4218, Q(179) 
                           => n_4219, Q(178) => n_4220, Q(177) => n_4221, 
                           Q(176) => n_4222, Q(175) => n_4223, Q(174) => n_4224
                           , Q(173) => n_4225, Q(172) => n_4226, Q(171) => 
                           n_4227, Q(170) => n_4228, Q(169) => n_4229, Q(168) 
                           => n_4230, Q(167) => n_4231, Q(166) => n_4232, 
                           Q(165) => n_4233, Q(164) => n_4234, Q(163) => n_4235
                           , Q(162) => n_4236, Q(161) => n_4237, Q(160) => 
                           n_4238, Q(159) => n_4239, Q(158) => n_4240, Q(157) 
                           => n_4241, Q(156) => n_4242, Q(155) => n_4243, 
                           Q(154) => n_4244, Q(153) => n_4245, Q(152) => n_4246
                           , Q(151) => n_4247, Q(150) => n_4248, Q(149) => 
                           n_4249, Q(148) => n_4250, Q(147) => n_4251, Q(146) 
                           => n_4252, Q(145) => n_4253, Q(144) => n_4254, 
                           Q(143) => n_4255, Q(142) => n_4256, Q(141) => n_4257
                           , Q(140) => n_4258, Q(139) => n_4259, Q(138) => 
                           n_4260, Q(137) => n_4261, Q(136) => n_4262, Q(135) 
                           => n_4263, Q(134) => n_4264, Q(133) => n_4265, 
                           Q(132) => n_4266, Q(131) => n_4267, Q(130) => n_4268
                           , Q(129) => n_4269, Q(128) => n_4270, Q(127) => 
                           n_4271, Q(126) => n_4272, Q(125) => n_4273, Q(124) 
                           => n_4274, Q(123) => n_4275, Q(122) => n_4276, 
                           Q(121) => n_4277, Q(120) => n_4278, Q(119) => n_4279
                           , Q(118) => n_4280, Q(117) => n_4281, Q(116) => 
                           n_4282, Q(115) => n_4283, Q(114) => n_4284, Q(113) 
                           => n_4285, Q(112) => n_4286, Q(111) => n_4287, 
                           Q(110) => n_4288, Q(109) => n_4289, Q(108) => n_4290
                           , Q(107) => n_4291, Q(106) => n_4292, Q(105) => 
                           n_4293, Q(104) => n_4294, Q(103) => n_4295, Q(102) 
                           => n_4296, Q(101) => n_4297, Q(100) => n_4298, Q(99)
                           => n_4299, Q(98) => n_4300, Q(97) => n_4301, Q(96) 
                           => n_4302, Q(95) => n_4303, Q(94) => n_4304, Q(93) 
                           => n_4305, Q(92) => n_4306, Q(91) => n_4307, Q(90) 
                           => n_4308, Q(89) => n_4309, Q(88) => n_4310, Q(87) 
                           => n_4311, Q(86) => n_4312, Q(85) => n_4313, Q(84) 
                           => n_4314, Q(83) => n_4315, Q(82) => n_4316, Q(81) 
                           => n_4317, Q(80) => n_4318, Q(79) => n_4319, Q(78) 
                           => n_4320, Q(77) => n_4321, Q(76) => n_4322, Q(75) 
                           => n_4323, Q(74) => n_4324, Q(73) => n_4325, Q(72) 
                           => n_4326, Q(71) => n_4327, Q(70) => n_4328, Q(69) 
                           => n_4329, Q(68) => n_4330, Q(67) => n_4331, Q(66) 
                           => n_4332, Q(65) => n_4333, Q(64) => n_4334, Q(63) 
                           => n_4335, Q(62) => n_4336, Q(61) => n_4337, Q(60) 
                           => n_4338, Q(59) => n_4339, Q(58) => n_4340, Q(57) 
                           => n_4341, Q(56) => n_4342, Q(55) => n_4343, Q(54) 
                           => n_4344, Q(53) => n_4345, Q(52) => n_4346, Q(51) 
                           => n_4347, Q(50) => n_4348, Q(49) => n_4349, Q(48) 
                           => n_4350, Q(47) => n_4351, Q(46) => n_4352, Q(45) 
                           => n_4353, Q(44) => n_4354, Q(43) => n_4355, Q(42) 
                           => n_4356, Q(41) => n_4357, Q(40) => n_4358, Q(39) 
                           => n_4359, Q(38) => n_4360, Q(37) => n_4361, Q(36) 
                           => n_4362, Q(35) => n_4363, Q(34) => n_4364, Q(33) 
                           => n_4365, Q(32) => n_4366, Q(31) => n_4367, Q(30) 
                           => n_4368, Q(29) => n_4369, Q(28) => n_4370, Q(27) 
                           => n_4371, Q(26) => n_4372, Q(25) => n_4373, Q(24) 
                           => n_4374, Q(23) => n_4375, Q(22) => n_4376, Q(21) 
                           => n_4377, Q(20) => n_4378, Q(19) => n_4379, Q(18) 
                           => n_4380, Q(17) => n_4381, Q(16) => n_4382, Q(15) 
                           => n_4383, Q(14) => n_4384, Q(13) => n_4385, Q(12) 
                           => n_4386, Q(11) => n_4387, Q(10) => n_4388, Q(9) =>
                           n_4389, Q(8) => n_4390, Q(7) => n_4391, Q(6) => 
                           n_4392, Q(5) => n_4393, Q(4) => n_4394, Q(3) => 
                           n_4395, Q(2) => n_4396, Q(1) => n_4397, Q(0) => 
                           n_4398);
   MUXi_7 : MUX_zbit_nbit_N31_Z3 port map( inputs(0) => X_Logic0_port, 
                           inputs(1) => X_Logic0_port, inputs(2) => 
                           X_Logic0_port, inputs(3) => X_Logic0_port, inputs(4)
                           => X_Logic0_port, inputs(5) => X_Logic0_port, 
                           inputs(6) => X_Logic0_port, inputs(7) => 
                           X_Logic0_port, inputs(8) => X_Logic0_port, inputs(9)
                           => X_Logic0_port, inputs(10) => X_Logic0_port, 
                           inputs(11) => X_Logic0_port, inputs(12) => 
                           X_Logic0_port, inputs(13) => X_Logic0_port, 
                           inputs(14) => X_Logic0_port, inputs(15) => 
                           X_Logic0_port, inputs(16) => X_Logic0_port, 
                           inputs(17) => X_Logic0_port, inputs(18) => 
                           X_Logic0_port, inputs(19) => X_Logic0_port, 
                           inputs(20) => X_Logic0_port, inputs(21) => 
                           X_Logic0_port, inputs(22) => X_Logic0_port, 
                           inputs(23) => X_Logic0_port, inputs(24) => 
                           X_Logic0_port, inputs(25) => X_Logic0_port, 
                           inputs(26) => X_Logic0_port, inputs(27) => 
                           X_Logic0_port, inputs(28) => X_Logic0_port, 
                           inputs(29) => X_Logic0_port, inputs(30) => 
                           X_Logic0_port, inputs(31) => muxes_in_7_31_port, 
                           inputs(32) => muxes_in_7_32_port, inputs(33) => 
                           muxes_in_7_33_port, inputs(34) => muxes_in_7_34_port
                           , inputs(35) => muxes_in_7_35_port, inputs(36) => 
                           muxes_in_7_36_port, inputs(37) => muxes_in_7_37_port
                           , inputs(38) => muxes_in_7_38_port, inputs(39) => 
                           muxes_in_7_39_port, inputs(40) => muxes_in_7_40_port
                           , inputs(41) => muxes_in_7_41_port, inputs(42) => 
                           muxes_in_7_42_port, inputs(43) => muxes_in_7_43_port
                           , inputs(44) => muxes_in_7_44_port, inputs(45) => 
                           muxes_in_7_45_port, inputs(46) => muxes_in_7_46_port
                           , inputs(47) => muxes_in_7_47_port, inputs(48) => 
                           muxes_in_7_48_port, inputs(49) => muxes_in_7_49_port
                           , inputs(50) => muxes_in_7_50_port, inputs(51) => 
                           muxes_in_7_51_port, inputs(52) => muxes_in_7_52_port
                           , inputs(53) => muxes_in_7_53_port, inputs(54) => 
                           muxes_in_7_54_port, inputs(55) => muxes_in_7_55_port
                           , inputs(56) => muxes_in_7_56_port, inputs(57) => 
                           muxes_in_7_57_port, inputs(58) => muxes_in_7_58_port
                           , inputs(59) => muxes_in_7_59_port, inputs(60) => 
                           X_Logic0_port, inputs(61) => X_Logic0_port, 
                           inputs(62) => muxes_in_7_62_port, inputs(63) => 
                           muxes_in_7_63_port, inputs(64) => muxes_in_7_64_port
                           , inputs(65) => muxes_in_7_65_port, inputs(66) => 
                           muxes_in_7_66_port, inputs(67) => muxes_in_7_67_port
                           , inputs(68) => muxes_in_7_68_port, inputs(69) => 
                           muxes_in_7_69_port, inputs(70) => muxes_in_7_70_port
                           , inputs(71) => muxes_in_7_71_port, inputs(72) => 
                           muxes_in_7_72_port, inputs(73) => muxes_in_7_73_port
                           , inputs(74) => muxes_in_7_74_port, inputs(75) => 
                           muxes_in_7_75_port, inputs(76) => muxes_in_7_76_port
                           , inputs(77) => muxes_in_7_77_port, inputs(78) => 
                           muxes_in_7_78_port, inputs(79) => muxes_in_7_79_port
                           , inputs(80) => muxes_in_7_80_port, inputs(81) => 
                           muxes_in_7_81_port, inputs(82) => muxes_in_7_82_port
                           , inputs(83) => muxes_in_7_83_port, inputs(84) => 
                           muxes_in_7_84_port, inputs(85) => muxes_in_7_85_port
                           , inputs(86) => muxes_in_7_86_port, inputs(87) => 
                           muxes_in_7_87_port, inputs(88) => muxes_in_7_88_port
                           , inputs(89) => muxes_in_7_89_port, inputs(90) => 
                           muxes_in_7_90_port, inputs(91) => X_Logic0_port, 
                           inputs(92) => X_Logic0_port, inputs(93) => 
                           X_Logic0_port, inputs(94) => X_Logic0_port, 
                           inputs(95) => X_Logic0_port, inputs(96) => 
                           X_Logic0_port, inputs(97) => X_Logic0_port, 
                           inputs(98) => X_Logic0_port, inputs(99) => 
                           X_Logic0_port, inputs(100) => X_Logic0_port, 
                           inputs(101) => X_Logic0_port, inputs(102) => 
                           X_Logic0_port, inputs(103) => X_Logic0_port, 
                           inputs(104) => X_Logic0_port, inputs(105) => 
                           X_Logic0_port, inputs(106) => X_Logic0_port, 
                           inputs(107) => X_Logic0_port, inputs(108) => 
                           X_Logic0_port, inputs(109) => X_Logic0_port, 
                           inputs(110) => X_Logic0_port, inputs(111) => 
                           X_Logic0_port, inputs(112) => X_Logic0_port, 
                           inputs(113) => X_Logic0_port, inputs(114) => 
                           X_Logic0_port, inputs(115) => X_Logic0_port, 
                           inputs(116) => X_Logic0_port, inputs(117) => 
                           X_Logic0_port, inputs(118) => X_Logic0_port, 
                           inputs(119) => X_Logic0_port, inputs(120) => 
                           X_Logic0_port, inputs(121) => X_Logic0_port, 
                           inputs(122) => X_Logic0_port, inputs(123) => 
                           X_Logic0_port, inputs(124) => X_Logic0_port, 
                           inputs(125) => X_Logic0_port, inputs(126) => 
                           X_Logic0_port, inputs(127) => X_Logic0_port, 
                           inputs(128) => X_Logic0_port, inputs(129) => 
                           X_Logic0_port, inputs(130) => X_Logic0_port, 
                           inputs(131) => X_Logic0_port, inputs(132) => 
                           X_Logic0_port, inputs(133) => X_Logic0_port, 
                           inputs(134) => X_Logic0_port, inputs(135) => 
                           X_Logic0_port, inputs(136) => X_Logic0_port, 
                           inputs(137) => X_Logic0_port, inputs(138) => 
                           X_Logic0_port, inputs(139) => X_Logic0_port, 
                           inputs(140) => X_Logic0_port, inputs(141) => 
                           X_Logic0_port, inputs(142) => X_Logic0_port, 
                           inputs(143) => X_Logic0_port, inputs(144) => 
                           X_Logic0_port, inputs(145) => X_Logic0_port, 
                           inputs(146) => X_Logic0_port, inputs(147) => 
                           X_Logic0_port, inputs(148) => X_Logic0_port, 
                           inputs(149) => X_Logic0_port, inputs(150) => 
                           X_Logic0_port, inputs(151) => X_Logic0_port, 
                           inputs(152) => X_Logic0_port, inputs(153) => 
                           X_Logic0_port, inputs(154) => X_Logic0_port, 
                           inputs(155) => X_Logic0_port, inputs(156) => 
                           X_Logic0_port, inputs(157) => X_Logic0_port, 
                           inputs(158) => X_Logic0_port, inputs(159) => 
                           X_Logic0_port, inputs(160) => X_Logic0_port, 
                           inputs(161) => X_Logic0_port, inputs(162) => 
                           X_Logic0_port, inputs(163) => X_Logic0_port, 
                           inputs(164) => X_Logic0_port, inputs(165) => 
                           X_Logic0_port, inputs(166) => X_Logic0_port, 
                           inputs(167) => X_Logic0_port, inputs(168) => 
                           X_Logic0_port, inputs(169) => X_Logic0_port, 
                           inputs(170) => X_Logic0_port, inputs(171) => 
                           X_Logic0_port, inputs(172) => X_Logic0_port, 
                           inputs(173) => X_Logic0_port, inputs(174) => 
                           X_Logic0_port, inputs(175) => X_Logic0_port, 
                           inputs(176) => X_Logic0_port, inputs(177) => 
                           X_Logic0_port, inputs(178) => X_Logic0_port, 
                           inputs(179) => X_Logic0_port, inputs(180) => 
                           X_Logic0_port, inputs(181) => X_Logic0_port, 
                           inputs(182) => X_Logic0_port, inputs(183) => 
                           X_Logic0_port, inputs(184) => X_Logic0_port, 
                           inputs(185) => X_Logic0_port, inputs(186) => 
                           muxes_in_7_186_port, inputs(187) => 
                           muxes_in_7_187_port, inputs(188) => 
                           muxes_in_7_188_port, inputs(189) => 
                           muxes_in_7_189_port, inputs(190) => 
                           muxes_in_7_190_port, inputs(191) => 
                           muxes_in_7_191_port, inputs(192) => 
                           muxes_in_7_192_port, inputs(193) => 
                           muxes_in_7_193_port, inputs(194) => 
                           muxes_in_7_194_port, inputs(195) => 
                           muxes_in_7_195_port, inputs(196) => 
                           muxes_in_7_196_port, inputs(197) => 
                           muxes_in_7_197_port, inputs(198) => 
                           muxes_in_7_198_port, inputs(199) => 
                           muxes_in_7_199_port, inputs(200) => 
                           muxes_in_7_200_port, inputs(201) => 
                           muxes_in_7_201_port, inputs(202) => 
                           muxes_in_7_202_port, inputs(203) => 
                           muxes_in_7_203_port, inputs(204) => 
                           muxes_in_7_204_port, inputs(205) => 
                           muxes_in_7_205_port, inputs(206) => 
                           muxes_in_7_206_port, inputs(207) => 
                           muxes_in_7_207_port, inputs(208) => 
                           muxes_in_7_208_port, inputs(209) => 
                           muxes_in_7_209_port, inputs(210) => 
                           muxes_in_7_210_port, inputs(211) => 
                           muxes_in_7_211_port, inputs(212) => 
                           muxes_in_7_212_port, inputs(213) => 
                           muxes_in_7_213_port, inputs(214) => 
                           muxes_in_7_214_port, inputs(215) => X_Logic0_port, 
                           inputs(216) => X_Logic0_port, inputs(217) => 
                           muxes_in_7_217_port, inputs(218) => 
                           muxes_in_7_218_port, inputs(219) => 
                           muxes_in_7_219_port, inputs(220) => 
                           muxes_in_7_220_port, inputs(221) => 
                           muxes_in_7_221_port, inputs(222) => 
                           muxes_in_7_222_port, inputs(223) => 
                           muxes_in_7_223_port, inputs(224) => 
                           muxes_in_7_224_port, inputs(225) => 
                           muxes_in_7_225_port, inputs(226) => 
                           muxes_in_7_226_port, inputs(227) => 
                           muxes_in_7_227_port, inputs(228) => 
                           muxes_in_7_228_port, inputs(229) => 
                           muxes_in_7_229_port, inputs(230) => 
                           muxes_in_7_230_port, inputs(231) => 
                           muxes_in_7_231_port, inputs(232) => 
                           muxes_in_7_232_port, inputs(233) => 
                           muxes_in_7_233_port, inputs(234) => 
                           muxes_in_7_234_port, inputs(235) => 
                           muxes_in_7_235_port, inputs(236) => 
                           muxes_in_7_236_port, inputs(237) => 
                           muxes_in_7_237_port, inputs(238) => 
                           muxes_in_7_238_port, inputs(239) => 
                           muxes_in_7_239_port, inputs(240) => 
                           muxes_in_7_240_port, inputs(241) => 
                           muxes_in_7_241_port, inputs(242) => 
                           muxes_in_7_242_port, inputs(243) => 
                           muxes_in_7_243_port, inputs(244) => 
                           muxes_in_7_244_port, inputs(245) => 
                           muxes_in_7_245_port, inputs(246) => X_Logic0_port, 
                           inputs(247) => X_Logic0_port, SEL(2) => 
                           encoder_out_7_2_port, SEL(1) => encoder_out_7_1_port
                           , SEL(0) => encoder_out_7_0_port, Y(30) => 
                           mux_out_7_30_port, Y(29) => mux_out_7_29_port, Y(28)
                           => mux_out_7_28_port, Y(27) => mux_out_7_27_port, 
                           Y(26) => mux_out_7_26_port, Y(25) => 
                           mux_out_7_25_port, Y(24) => mux_out_7_24_port, Y(23)
                           => mux_out_7_23_port, Y(22) => mux_out_7_22_port, 
                           Y(21) => mux_out_7_21_port, Y(20) => 
                           mux_out_7_20_port, Y(19) => mux_out_7_19_port, Y(18)
                           => mux_out_7_18_port, Y(17) => mux_out_7_17_port, 
                           Y(16) => mux_out_7_16_port, Y(15) => 
                           mux_out_7_15_port, Y(14) => mux_out_7_14_port, Y(13)
                           => mux_out_7_13_port, Y(12) => mux_out_7_12_port, 
                           Y(11) => mux_out_7_11_port, Y(10) => 
                           mux_out_7_10_port, Y(9) => mux_out_7_9_port, Y(8) =>
                           mux_out_7_8_port, Y(7) => mux_out_7_7_port, Y(6) => 
                           mux_out_7_6_port, Y(5) => mux_out_7_5_port, Y(4) => 
                           mux_out_7_4_port, Y(3) => mux_out_7_3_port, Y(2) => 
                           mux_out_7_2_port, Y(1) => mux_out_7_1_port, Y(0) => 
                           mux_out_7_0_port);
   ADDn_7 : adder_NBIT31 port map( a(30) => mux_out_7_30_port, a(29) => 
                           mux_out_7_29_port, a(28) => mux_out_7_28_port, a(27)
                           => mux_out_7_27_port, a(26) => mux_out_7_26_port, 
                           a(25) => mux_out_7_25_port, a(24) => 
                           mux_out_7_24_port, a(23) => mux_out_7_23_port, a(22)
                           => mux_out_7_22_port, a(21) => mux_out_7_21_port, 
                           a(20) => mux_out_7_20_port, a(19) => 
                           mux_out_7_19_port, a(18) => mux_out_7_18_port, a(17)
                           => mux_out_7_17_port, a(16) => mux_out_7_16_port, 
                           a(15) => mux_out_7_15_port, a(14) => 
                           mux_out_7_14_port, a(13) => mux_out_7_13_port, a(12)
                           => mux_out_7_12_port, a(11) => mux_out_7_11_port, 
                           a(10) => mux_out_7_10_port, a(9) => mux_out_7_9_port
                           , a(8) => mux_out_7_8_port, a(7) => mux_out_7_7_port
                           , a(6) => mux_out_7_6_port, a(5) => mux_out_7_5_port
                           , a(4) => mux_out_7_4_port, a(3) => mux_out_7_3_port
                           , a(2) => mux_out_7_2_port, a(1) => mux_out_7_1_port
                           , a(0) => mux_out_7_0_port, b(30) => 
                           sum_B_in_7_30_port, b(29) => sum_B_in_7_30_port, 
                           b(28) => sum_B_in_7_30_port, b(27) => 
                           sum_B_in_7_27_port, b(26) => sum_B_in_7_26_port, 
                           b(25) => sum_B_in_7_25_port, b(24) => 
                           sum_B_in_7_24_port, b(23) => sum_B_in_7_23_port, 
                           b(22) => sum_B_in_7_22_port, b(21) => 
                           sum_B_in_7_21_port, b(20) => sum_B_in_7_20_port, 
                           b(19) => sum_B_in_7_19_port, b(18) => 
                           sum_B_in_7_18_port, b(17) => sum_B_in_7_17_port, 
                           b(16) => sum_B_in_7_16_port, b(15) => 
                           sum_B_in_7_15_port, b(14) => sum_B_in_7_14_port, 
                           b(13) => sum_B_in_7_13_port, b(12) => 
                           sum_B_in_7_12_port, b(11) => sum_B_in_7_11_port, 
                           b(10) => sum_B_in_7_10_port, b(9) => 
                           sum_B_in_7_9_port, b(8) => sum_B_in_7_8_port, b(7) 
                           => sum_B_in_7_7_port, b(6) => sum_B_in_7_6_port, 
                           b(5) => sum_B_in_7_5_port, b(4) => sum_B_in_7_4_port
                           , b(3) => sum_B_in_7_3_port, b(2) => 
                           sum_B_in_7_2_port, b(1) => sum_B_in_7_1_port, b(0) 
                           => sum_B_in_7_0_port, cin => X_Logic0_port, s(31) =>
                           result(31), s(30) => result(30), s(29) => result(29)
                           , s(28) => result(28), s(27) => result(27), s(26) =>
                           result(26), s(25) => result(25), s(24) => result(24)
                           , s(23) => result(23), s(22) => result(22), s(21) =>
                           result(21), s(20) => result(20), s(19) => result(19)
                           , s(18) => result(18), s(17) => result(17), s(16) =>
                           result(16), s(15) => result(15), s(14) => result(14)
                           , s(13) => result(13), s(12) => result(12), s(11) =>
                           result(11), s(10) => result(10), s(9) => result(9), 
                           s(8) => result(8), s(7) => result(7), s(6) => 
                           result(6), s(5) => result(5), s(4) => result(4), 
                           s(3) => result(3), s(2) => result(2), s(1) => 
                           result(1), s(0) => result(0));
   pip_del_reg_i_2 : reg_nbit_n16_0 port map( clk => n11, reset => n4, d(15) =>
                           multiplicand(15), d(14) => multiplicand(14), d(13) 
                           => multiplicand(13), d(12) => multiplicand(12), 
                           d(11) => multiplicand(11), d(10) => multiplicand(10)
                           , d(9) => multiplicand(9), d(8) => multiplicand(8), 
                           d(7) => multiplicand(7), d(6) => multiplicand(6), 
                           d(5) => multiplicand(5), d(4) => multiplicand(4), 
                           d(3) => multiplicand(3), d(2) => multiplicand(2), 
                           d(1) => multiplicand(1), d(0) => multiplicand(0), 
                           Q(15) => multiplicand_pip_2_15_port, Q(14) => 
                           multiplicand_pip_2_14_port, Q(13) => 
                           multiplicand_pip_2_13_port, Q(12) => 
                           multiplicand_pip_2_12_port, Q(11) => 
                           multiplicand_pip_2_11_port, Q(10) => 
                           multiplicand_pip_2_10_port, Q(9) => 
                           multiplicand_pip_2_9_port, Q(8) => 
                           multiplicand_pip_2_8_port, Q(7) => 
                           multiplicand_pip_2_7_port, Q(6) => 
                           multiplicand_pip_2_6_port, Q(5) => 
                           multiplicand_pip_2_5_port, Q(4) => 
                           multiplicand_pip_2_4_port, Q(3) => 
                           multiplicand_pip_2_3_port, Q(2) => 
                           multiplicand_pip_2_2_port, Q(1) => 
                           multiplicand_pip_2_1_port, Q(0) => 
                           multiplicand_pip_2_0_port);
   pip_del_reg_i_3 : reg_nbit_n16_5 port map( clk => n11, reset => n3, d(15) =>
                           multiplicand_pip_2_15_port, d(14) => 
                           multiplicand_pip_2_14_port, d(13) => 
                           multiplicand_pip_2_13_port, d(12) => 
                           multiplicand_pip_2_12_port, d(11) => 
                           multiplicand_pip_2_11_port, d(10) => 
                           multiplicand_pip_2_10_port, d(9) => 
                           multiplicand_pip_2_9_port, d(8) => 
                           multiplicand_pip_2_8_port, d(7) => 
                           multiplicand_pip_2_7_port, d(6) => 
                           multiplicand_pip_2_6_port, d(5) => 
                           multiplicand_pip_2_5_port, d(4) => 
                           multiplicand_pip_2_4_port, d(3) => 
                           multiplicand_pip_2_3_port, d(2) => 
                           multiplicand_pip_2_2_port, d(1) => 
                           multiplicand_pip_2_1_port, d(0) => 
                           multiplicand_pip_2_0_port, Q(15) => 
                           multiplicand_pip_3_15_port, Q(14) => 
                           multiplicand_pip_3_14_port, Q(13) => 
                           multiplicand_pip_3_13_port, Q(12) => 
                           multiplicand_pip_3_12_port, Q(11) => 
                           multiplicand_pip_3_11_port, Q(10) => 
                           multiplicand_pip_3_10_port, Q(9) => 
                           multiplicand_pip_3_9_port, Q(8) => 
                           multiplicand_pip_3_8_port, Q(7) => 
                           multiplicand_pip_3_7_port, Q(6) => 
                           multiplicand_pip_3_6_port, Q(5) => 
                           multiplicand_pip_3_5_port, Q(4) => 
                           multiplicand_pip_3_4_port, Q(3) => 
                           multiplicand_pip_3_3_port, Q(2) => 
                           multiplicand_pip_3_2_port, Q(1) => 
                           multiplicand_pip_3_1_port, Q(0) => 
                           multiplicand_pip_3_0_port);
   pip_del_reg_i_4 : reg_nbit_n16_4 port map( clk => n11, reset => n3, d(15) =>
                           multiplicand_pip_3_15_port, d(14) => 
                           multiplicand_pip_3_14_port, d(13) => 
                           multiplicand_pip_3_13_port, d(12) => 
                           multiplicand_pip_3_12_port, d(11) => 
                           multiplicand_pip_3_11_port, d(10) => 
                           multiplicand_pip_3_10_port, d(9) => 
                           multiplicand_pip_3_9_port, d(8) => 
                           multiplicand_pip_3_8_port, d(7) => 
                           multiplicand_pip_3_7_port, d(6) => 
                           multiplicand_pip_3_6_port, d(5) => 
                           multiplicand_pip_3_5_port, d(4) => 
                           multiplicand_pip_3_4_port, d(3) => 
                           multiplicand_pip_3_3_port, d(2) => 
                           multiplicand_pip_3_2_port, d(1) => 
                           multiplicand_pip_3_1_port, d(0) => 
                           multiplicand_pip_3_0_port, Q(15) => 
                           multiplicand_pip_4_15_port, Q(14) => 
                           multiplicand_pip_4_14_port, Q(13) => 
                           multiplicand_pip_4_13_port, Q(12) => 
                           multiplicand_pip_4_12_port, Q(11) => 
                           multiplicand_pip_4_11_port, Q(10) => 
                           multiplicand_pip_4_10_port, Q(9) => 
                           multiplicand_pip_4_9_port, Q(8) => 
                           multiplicand_pip_4_8_port, Q(7) => 
                           multiplicand_pip_4_7_port, Q(6) => 
                           multiplicand_pip_4_6_port, Q(5) => 
                           multiplicand_pip_4_5_port, Q(4) => 
                           multiplicand_pip_4_4_port, Q(3) => 
                           multiplicand_pip_4_3_port, Q(2) => 
                           multiplicand_pip_4_2_port, Q(1) => 
                           multiplicand_pip_4_1_port, Q(0) => 
                           multiplicand_pip_4_0_port);
   pip_del_reg_i_5 : reg_nbit_n16_3 port map( clk => n12, reset => n3, d(15) =>
                           multiplicand_pip_4_15_port, d(14) => 
                           multiplicand_pip_4_14_port, d(13) => 
                           multiplicand_pip_4_13_port, d(12) => 
                           multiplicand_pip_4_12_port, d(11) => 
                           multiplicand_pip_4_11_port, d(10) => 
                           multiplicand_pip_4_10_port, d(9) => 
                           multiplicand_pip_4_9_port, d(8) => 
                           multiplicand_pip_4_8_port, d(7) => 
                           multiplicand_pip_4_7_port, d(6) => 
                           multiplicand_pip_4_6_port, d(5) => 
                           multiplicand_pip_4_5_port, d(4) => 
                           multiplicand_pip_4_4_port, d(3) => 
                           multiplicand_pip_4_3_port, d(2) => 
                           multiplicand_pip_4_2_port, d(1) => 
                           multiplicand_pip_4_1_port, d(0) => 
                           multiplicand_pip_4_0_port, Q(15) => 
                           multiplicand_pip_5_15_port, Q(14) => 
                           multiplicand_pip_5_14_port, Q(13) => 
                           multiplicand_pip_5_13_port, Q(12) => 
                           multiplicand_pip_5_12_port, Q(11) => 
                           multiplicand_pip_5_11_port, Q(10) => 
                           multiplicand_pip_5_10_port, Q(9) => 
                           multiplicand_pip_5_9_port, Q(8) => 
                           multiplicand_pip_5_8_port, Q(7) => 
                           multiplicand_pip_5_7_port, Q(6) => 
                           multiplicand_pip_5_6_port, Q(5) => 
                           multiplicand_pip_5_5_port, Q(4) => 
                           multiplicand_pip_5_4_port, Q(3) => 
                           multiplicand_pip_5_3_port, Q(2) => 
                           multiplicand_pip_5_2_port, Q(1) => 
                           multiplicand_pip_5_1_port, Q(0) => 
                           multiplicand_pip_5_0_port);
   pip_del_reg_i_6 : reg_nbit_n16_2 port map( clk => n12, reset => n4, d(15) =>
                           multiplicand_pip_5_15_port, d(14) => 
                           multiplicand_pip_5_14_port, d(13) => 
                           multiplicand_pip_5_13_port, d(12) => 
                           multiplicand_pip_5_12_port, d(11) => 
                           multiplicand_pip_5_11_port, d(10) => 
                           multiplicand_pip_5_10_port, d(9) => 
                           multiplicand_pip_5_9_port, d(8) => 
                           multiplicand_pip_5_8_port, d(7) => 
                           multiplicand_pip_5_7_port, d(6) => 
                           multiplicand_pip_5_6_port, d(5) => 
                           multiplicand_pip_5_5_port, d(4) => 
                           multiplicand_pip_5_4_port, d(3) => 
                           multiplicand_pip_5_3_port, d(2) => 
                           multiplicand_pip_5_2_port, d(1) => 
                           multiplicand_pip_5_1_port, d(0) => 
                           multiplicand_pip_5_0_port, Q(15) => 
                           multiplicand_pip_6_15_port, Q(14) => 
                           multiplicand_pip_6_14_port, Q(13) => 
                           multiplicand_pip_6_13_port, Q(12) => 
                           multiplicand_pip_6_12_port, Q(11) => 
                           multiplicand_pip_6_11_port, Q(10) => 
                           multiplicand_pip_6_10_port, Q(9) => 
                           multiplicand_pip_6_9_port, Q(8) => 
                           multiplicand_pip_6_8_port, Q(7) => 
                           multiplicand_pip_6_7_port, Q(6) => 
                           multiplicand_pip_6_6_port, Q(5) => 
                           multiplicand_pip_6_5_port, Q(4) => 
                           multiplicand_pip_6_4_port, Q(3) => 
                           multiplicand_pip_6_3_port, Q(2) => 
                           multiplicand_pip_6_2_port, Q(1) => 
                           multiplicand_pip_6_1_port, Q(0) => 
                           multiplicand_pip_6_0_port);
   pip_del_reg_i_7 : reg_nbit_n16_1 port map( clk => n11, reset => n4, d(15) =>
                           multiplicand_pip_6_15_port, d(14) => 
                           multiplicand_pip_6_14_port, d(13) => 
                           multiplicand_pip_6_13_port, d(12) => 
                           multiplicand_pip_6_12_port, d(11) => 
                           multiplicand_pip_6_11_port, d(10) => 
                           multiplicand_pip_6_10_port, d(9) => 
                           multiplicand_pip_6_9_port, d(8) => 
                           multiplicand_pip_6_8_port, d(7) => 
                           multiplicand_pip_6_7_port, d(6) => 
                           multiplicand_pip_6_6_port, d(5) => 
                           multiplicand_pip_6_5_port, d(4) => 
                           multiplicand_pip_6_4_port, d(3) => 
                           multiplicand_pip_6_3_port, d(2) => 
                           multiplicand_pip_6_2_port, d(1) => 
                           multiplicand_pip_6_1_port, d(0) => 
                           multiplicand_pip_6_0_port, Q(15) => 
                           multiplicand_pip_7_15_port, Q(14) => 
                           multiplicand_pip_7_14_port, Q(13) => 
                           multiplicand_pip_7_13_port, Q(12) => n_4399, Q(11) 
                           => n_4400, Q(10) => n_4401, Q(9) => n_4402, Q(8) => 
                           n_4403, Q(7) => n_4404, Q(6) => n_4405, Q(5) => 
                           n_4406, Q(4) => n_4407, Q(3) => n_4408, Q(2) => 
                           n_4409, Q(1) => n_4410, Q(0) => n_4411);
   U2 : BUF_X1 port map( A => n2, Z => n5);
   U3 : BUF_X1 port map( A => n2, Z => n6);
   U4 : BUF_X1 port map( A => n1, Z => n3);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n8, Z => n12);
   U7 : BUF_X1 port map( A => n8, Z => n11);
   U8 : BUF_X1 port map( A => n7, Z => n10);
   U9 : BUF_X1 port map( A => n7, Z => n9);
   U10 : BUF_X1 port map( A => rst, Z => n2);
   U11 : BUF_X1 port map( A => rst, Z => n1);
   U12 : BUF_X1 port map( A => clk, Z => n7);
   U13 : BUF_X1 port map( A => clk, Z => n8);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity p4_adder_NBIT32 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end p4_adder_NBIT32;

architecture SYN_struc of p4_adder_NBIT32 is

   component SUM_GEN_NBIT32_NBLOCKS4
      port( A, B, Ci : in std_logic_vector (31 downto 0);  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component STCG_NBIT32_SDIST4
      port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            Cout : out std_logic_vector (32 downto 0));
   end component;
   
   signal C_select_31_port, C_select_30_port, C_select_29_port, 
      C_select_28_port, C_select_27_port, C_select_26_port, C_select_25_port, 
      C_select_24_port, C_select_23_port, C_select_22_port, C_select_21_port, 
      C_select_20_port, C_select_19_port, C_select_18_port, C_select_17_port, 
      C_select_16_port, C_select_15_port, C_select_14_port, C_select_13_port, 
      C_select_12_port, C_select_11_port, C_select_10_port, C_select_9_port, 
      C_select_8_port, C_select_7_port, C_select_6_port, C_select_5_port, 
      C_select_4_port, C_select_3_port, C_select_2_port, C_select_1_port, 
      C_select_0_port, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, 
      n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, 
      n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435 : 
      std_logic;

begin
   
   carry_select : STCG_NBIT32_SDIST4 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), B(31) => b(31), B(30) => b(30), 
                           B(29) => b(29), B(28) => b(28), B(27) => b(27), 
                           B(26) => b(26), B(25) => b(25), B(24) => b(24), 
                           B(23) => b(23), B(22) => b(22), B(21) => b(21), 
                           B(20) => b(20), B(19) => b(19), B(18) => b(18), 
                           B(17) => b(17), B(16) => b(16), B(15) => b(15), 
                           B(14) => b(14), B(13) => b(13), B(12) => b(12), 
                           B(11) => b(11), B(10) => b(10), B(9) => b(9), B(8) 
                           => b(8), B(7) => b(7), B(6) => b(6), B(5) => b(5), 
                           B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1) => 
                           b(1), B(0) => b(0), cin => cin, Cout(32) => cout, 
                           Cout(31) => n_4412, Cout(30) => n_4413, Cout(29) => 
                           n_4414, Cout(28) => C_select_28_port, Cout(27) => 
                           n_4415, Cout(26) => n_4416, Cout(25) => n_4417, 
                           Cout(24) => C_select_24_port, Cout(23) => n_4418, 
                           Cout(22) => n_4419, Cout(21) => n_4420, Cout(20) => 
                           C_select_20_port, Cout(19) => n_4421, Cout(18) => 
                           n_4422, Cout(17) => n_4423, Cout(16) => 
                           C_select_16_port, Cout(15) => n_4424, Cout(14) => 
                           n_4425, Cout(13) => n_4426, Cout(12) => 
                           C_select_12_port, Cout(11) => n_4427, Cout(10) => 
                           n_4428, Cout(9) => n_4429, Cout(8) => 
                           C_select_8_port, Cout(7) => n_4430, Cout(6) => 
                           n_4431, Cout(5) => n_4432, Cout(4) => 
                           C_select_4_port, Cout(3) => n_4433, Cout(2) => 
                           n_4434, Cout(1) => n_4435, Cout(0) => 
                           C_select_0_port);
   sums : SUM_GEN_NBIT32_NBLOCKS4 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), B(31) => b(31), B(30) => b(30), 
                           B(29) => b(29), B(28) => b(28), B(27) => b(27), 
                           B(26) => b(26), B(25) => b(25), B(24) => b(24), 
                           B(23) => b(23), B(22) => b(22), B(21) => b(21), 
                           B(20) => b(20), B(19) => b(19), B(18) => b(18), 
                           B(17) => b(17), B(16) => b(16), B(15) => b(15), 
                           B(14) => b(14), B(13) => b(13), B(12) => b(12), 
                           B(11) => b(11), B(10) => b(10), B(9) => b(9), B(8) 
                           => b(8), B(7) => b(7), B(6) => b(6), B(5) => b(5), 
                           B(4) => b(4), B(3) => b(3), B(2) => b(2), B(1) => 
                           b(1), B(0) => b(0), Ci(31) => C_select_31_port, 
                           Ci(30) => C_select_30_port, Ci(29) => 
                           C_select_29_port, Ci(28) => C_select_28_port, Ci(27)
                           => C_select_27_port, Ci(26) => C_select_26_port, 
                           Ci(25) => C_select_25_port, Ci(24) => 
                           C_select_24_port, Ci(23) => C_select_23_port, Ci(22)
                           => C_select_22_port, Ci(21) => C_select_21_port, 
                           Ci(20) => C_select_20_port, Ci(19) => 
                           C_select_19_port, Ci(18) => C_select_18_port, Ci(17)
                           => C_select_17_port, Ci(16) => C_select_16_port, 
                           Ci(15) => C_select_15_port, Ci(14) => 
                           C_select_14_port, Ci(13) => C_select_13_port, Ci(12)
                           => C_select_12_port, Ci(11) => C_select_11_port, 
                           Ci(10) => C_select_10_port, Ci(9) => C_select_9_port
                           , Ci(8) => C_select_8_port, Ci(7) => C_select_7_port
                           , Ci(6) => C_select_6_port, Ci(5) => C_select_5_port
                           , Ci(4) => C_select_4_port, Ci(3) => C_select_3_port
                           , Ci(2) => C_select_2_port, Ci(1) => C_select_1_port
                           , Ci(0) => C_select_0_port, S(31) => s(31), S(30) =>
                           s(30), S(29) => s(29), S(28) => s(28), S(27) => 
                           s(27), S(26) => s(26), S(25) => s(25), S(24) => 
                           s(24), S(23) => s(23), S(22) => s(22), S(21) => 
                           s(21), S(20) => s(20), S(19) => s(19), S(18) => 
                           s(18), S(17) => s(17), S(16) => s(16), S(15) => 
                           s(15), S(14) => s(14), S(13) => s(13), S(12) => 
                           s(12), S(11) => s(11), S(10) => s(10), S(9) => s(9),
                           S(8) => s(8), S(7) => s(7), S(6) => s(6), S(5) => 
                           s(5), S(4) => s(4), S(3) => s(3), S(2) => s(2), S(1)
                           => s(1), S(0) => s(0));
   C_select_1_port <= '0';
   C_select_2_port <= '0';
   C_select_3_port <= '0';
   C_select_5_port <= '0';
   C_select_6_port <= '0';
   C_select_7_port <= '0';
   C_select_9_port <= '0';
   C_select_10_port <= '0';
   C_select_11_port <= '0';
   C_select_13_port <= '0';
   C_select_14_port <= '0';
   C_select_15_port <= '0';
   C_select_17_port <= '0';
   C_select_18_port <= '0';
   C_select_19_port <= '0';
   C_select_21_port <= '0';
   C_select_22_port <= '0';
   C_select_23_port <= '0';
   C_select_25_port <= '0';
   C_select_26_port <= '0';
   C_select_27_port <= '0';
   C_select_29_port <= '0';
   C_select_30_port <= '0';
   C_select_31_port <= '0';

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk, rst : in std_logic;  zero_mul_detect, mul_exeception : out 
         std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         );

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component general_alu_N32_DW01_cmp6_1
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component general_alu_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component boothmul_pipelined_N16
      port( clk, rst : in std_logic;  multiplier, multiplicand : in 
            std_logic_vector (15 downto 0);  result : out std_logic_vector (31 
            downto 0));
   end component;
   
   component p4_adder_NBIT32
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      adder_out_31_port, adder_out_30_port, adder_out_29_port, 
      adder_out_28_port, adder_out_27_port, adder_out_26_port, 
      adder_out_25_port, adder_out_24_port, adder_out_23_port, 
      adder_out_22_port, adder_out_21_port, adder_out_20_port, 
      adder_out_19_port, adder_out_18_port, adder_out_17_port, 
      adder_out_16_port, adder_out_15_port, adder_out_14_port, 
      adder_out_13_port, adder_out_12_port, adder_out_11_port, 
      adder_out_10_port, adder_out_9_port, adder_out_8_port, adder_out_7_port, 
      adder_out_6_port, adder_out_5_port, adder_out_4_port, adder_out_3_port, 
      adder_out_2_port, adder_out_1_port, adder_out_0_port, cout, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, data2_mul_0_port, dataout_mul_31_port, 
      dataout_mul_30_port, dataout_mul_29_port, dataout_mul_28_port, 
      dataout_mul_27_port, dataout_mul_26_port, dataout_mul_25_port, 
      dataout_mul_24_port, dataout_mul_23_port, dataout_mul_22_port, 
      dataout_mul_21_port, dataout_mul_20_port, dataout_mul_19_port, 
      dataout_mul_18_port, dataout_mul_17_port, dataout_mul_16_port, 
      dataout_mul_15_port, dataout_mul_14_port, dataout_mul_13_port, 
      dataout_mul_12_port, dataout_mul_11_port, dataout_mul_10_port, 
      dataout_mul_9_port, dataout_mul_8_port, dataout_mul_7_port, 
      dataout_mul_6_port, dataout_mul_5_port, dataout_mul_4_port, 
      dataout_mul_3_port, dataout_mul_2_port, dataout_mul_1_port, 
      dataout_mul_0_port, check_mul_logic, N2513, N2514, N2515, N2517, N2518, 
      N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, 
      N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, 
      N2539, N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, n1,
      n98, n553, n554, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
      n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, 
      n_4444 : std_logic;

begin
   
   n1 <= '0';
   n98 <= '1';
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n554, Q => 
                           DATA2_I_31_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n554, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n554, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n554, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n554, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n554, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n554, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n554, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n554, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n554, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n554, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n554, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           data2_mul_0_port);
   check_mul_logic_reg : DLL_X1 port map( D => n1034, GN => n553, Q => 
                           check_mul_logic);
   p4_adder_lab : p4_adder_NBIT32 port map( a(31) => DATA1(31), a(30) => 
                           DATA1(30), a(29) => DATA1(29), a(28) => DATA1(28), 
                           a(27) => DATA1(27), a(26) => DATA1(26), a(25) => 
                           DATA1(25), a(24) => DATA1(24), a(23) => DATA1(23), 
                           a(22) => DATA1(22), a(21) => DATA1(21), a(20) => 
                           DATA1(20), a(19) => DATA1(19), a(18) => DATA1(18), 
                           a(17) => DATA1(17), a(16) => DATA1(16), a(15) => 
                           DATA1(15), a(14) => DATA1(14), a(13) => DATA1(13), 
                           a(12) => DATA1(12), a(11) => DATA1(11), a(10) => 
                           DATA1(10), a(9) => DATA1(9), a(8) => DATA1(8), a(7) 
                           => DATA1(7), a(6) => DATA1(6), a(5) => DATA1(5), 
                           a(4) => DATA1(4), a(3) => DATA1(3), a(2) => DATA1(2)
                           , a(1) => DATA1(1), a(0) => DATA1(0), b(31) => 
                           DATA2_I_31_port, b(30) => DATA2_I_30_port, b(29) => 
                           DATA2_I_29_port, b(28) => DATA2_I_28_port, b(27) => 
                           DATA2_I_27_port, b(26) => DATA2_I_26_port, b(25) => 
                           DATA2_I_25_port, b(24) => DATA2_I_24_port, b(23) => 
                           DATA2_I_23_port, b(22) => DATA2_I_22_port, b(21) => 
                           DATA2_I_21_port, b(20) => DATA2_I_20_port, b(19) => 
                           DATA2_I_19_port, b(18) => DATA2_I_18_port, b(17) => 
                           DATA2_I_17_port, b(16) => DATA2_I_16_port, b(15) => 
                           DATA2_I_15_port, b(14) => DATA2_I_14_port, b(13) => 
                           DATA2_I_13_port, b(12) => DATA2_I_12_port, b(11) => 
                           DATA2_I_11_port, b(10) => DATA2_I_10_port, b(9) => 
                           DATA2_I_9_port, b(8) => DATA2_I_8_port, b(7) => 
                           DATA2_I_7_port, b(6) => DATA2_I_6_port, b(5) => 
                           DATA2_I_5_port, b(4) => DATA2_I_4_port, b(3) => 
                           DATA2_I_3_port, b(2) => DATA2_I_2_port, b(1) => 
                           DATA2_I_1_port, b(0) => DATA2_I_0_port, cin => cin, 
                           s(31) => adder_out_31_port, s(30) => 
                           adder_out_30_port, s(29) => adder_out_29_port, s(28)
                           => adder_out_28_port, s(27) => adder_out_27_port, 
                           s(26) => adder_out_26_port, s(25) => 
                           adder_out_25_port, s(24) => adder_out_24_port, s(23)
                           => adder_out_23_port, s(22) => adder_out_22_port, 
                           s(21) => adder_out_21_port, s(20) => 
                           adder_out_20_port, s(19) => adder_out_19_port, s(18)
                           => adder_out_18_port, s(17) => adder_out_17_port, 
                           s(16) => adder_out_16_port, s(15) => 
                           adder_out_15_port, s(14) => adder_out_14_port, s(13)
                           => adder_out_13_port, s(12) => adder_out_12_port, 
                           s(11) => adder_out_11_port, s(10) => 
                           adder_out_10_port, s(9) => adder_out_9_port, s(8) =>
                           adder_out_8_port, s(7) => adder_out_7_port, s(6) => 
                           adder_out_6_port, s(5) => adder_out_5_port, s(4) => 
                           adder_out_4_port, s(3) => adder_out_3_port, s(2) => 
                           adder_out_2_port, s(1) => adder_out_1_port, s(0) => 
                           adder_out_0_port, cout => cout);
   boothmul_pipelined_i : boothmul_pipelined_N16 port map( clk => clk, rst => 
                           rst, multiplier(15) => data1_mul_15_port, 
                           multiplier(14) => data1_mul_14_port, multiplier(13) 
                           => data1_mul_13_port, multiplier(12) => 
                           data1_mul_12_port, multiplier(11) => 
                           data1_mul_11_port, multiplier(10) => 
                           data1_mul_10_port, multiplier(9) => data1_mul_9_port
                           , multiplier(8) => data1_mul_8_port, multiplier(7) 
                           => data1_mul_7_port, multiplier(6) => 
                           data1_mul_6_port, multiplier(5) => data1_mul_5_port,
                           multiplier(4) => data1_mul_4_port, multiplier(3) => 
                           data1_mul_3_port, multiplier(2) => data1_mul_2_port,
                           multiplier(1) => data1_mul_1_port, multiplier(0) => 
                           data1_mul_0_port, multiplicand(15) => 
                           data2_mul_15_port, multiplicand(14) => 
                           data2_mul_14_port, multiplicand(13) => 
                           data2_mul_13_port, multiplicand(12) => 
                           data2_mul_12_port, multiplicand(11) => 
                           data2_mul_11_port, multiplicand(10) => 
                           data2_mul_10_port, multiplicand(9) => 
                           data2_mul_9_port, multiplicand(8) => 
                           data2_mul_8_port, multiplicand(7) => 
                           data2_mul_7_port, multiplicand(6) => 
                           data2_mul_6_port, multiplicand(5) => 
                           data2_mul_5_port, multiplicand(4) => 
                           data2_mul_4_port, multiplicand(3) => 
                           data2_mul_3_port, multiplicand(2) => 
                           data2_mul_2_port, multiplicand(1) => 
                           data2_mul_1_port, multiplicand(0) => 
                           data2_mul_0_port, result(31) => dataout_mul_31_port,
                           result(30) => dataout_mul_30_port, result(29) => 
                           dataout_mul_29_port, result(28) => 
                           dataout_mul_28_port, result(27) => 
                           dataout_mul_27_port, result(26) => 
                           dataout_mul_26_port, result(25) => 
                           dataout_mul_25_port, result(24) => 
                           dataout_mul_24_port, result(23) => 
                           dataout_mul_23_port, result(22) => 
                           dataout_mul_22_port, result(21) => 
                           dataout_mul_21_port, result(20) => 
                           dataout_mul_20_port, result(19) => 
                           dataout_mul_19_port, result(18) => 
                           dataout_mul_18_port, result(17) => 
                           dataout_mul_17_port, result(16) => 
                           dataout_mul_16_port, result(15) => 
                           dataout_mul_15_port, result(14) => 
                           dataout_mul_14_port, result(13) => 
                           dataout_mul_13_port, result(12) => 
                           dataout_mul_12_port, result(11) => 
                           dataout_mul_11_port, result(10) => 
                           dataout_mul_10_port, result(9) => dataout_mul_9_port
                           , result(8) => dataout_mul_8_port, result(7) => 
                           dataout_mul_7_port, result(6) => dataout_mul_6_port,
                           result(5) => dataout_mul_5_port, result(4) => 
                           dataout_mul_4_port, result(3) => dataout_mul_3_port,
                           result(2) => dataout_mul_2_port, result(1) => 
                           dataout_mul_1_port, result(0) => dataout_mul_0_port)
                           ;
   ne_191 : general_alu_N32_DW01_cmp6_0 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(31) => 
                           DATA2(31), B(30) => DATA2(30), B(29) => DATA2(29), 
                           B(28) => DATA2(28), B(27) => DATA2(27), B(26) => 
                           DATA2(26), B(25) => DATA2(25), B(24) => DATA2(24), 
                           B(23) => DATA2(23), B(22) => DATA2(22), B(21) => 
                           DATA2(21), B(20) => DATA2(20), B(19) => DATA2(19), 
                           B(18) => DATA2(18), B(17) => DATA2(17), B(16) => 
                           DATA2(16), B(15) => DATA2(15), B(14) => DATA2(14), 
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), TC => n1, LT => n_4436, GT => n_4437, 
                           EQ => n_4438, LE => n_4439, GE => n_4440, NE => 
                           N2515);
   r323 : general_alu_N32_DW01_cmp6_1 port map( A(31) => DATA2(31), A(30) => 
                           DATA2(30), A(29) => DATA2(29), A(28) => DATA2(28), 
                           A(27) => DATA2(27), A(26) => DATA2(26), A(25) => 
                           DATA2(25), A(24) => DATA2(24), A(23) => DATA2(23), 
                           A(22) => DATA2(22), A(21) => DATA2(21), A(20) => 
                           DATA2(20), A(19) => DATA2(19), A(18) => DATA2(18), 
                           A(17) => DATA2(17), A(16) => DATA2(16), A(15) => 
                           DATA2(15), A(14) => DATA2(14), A(13) => DATA2(13), 
                           A(12) => DATA2(12), A(11) => DATA2(11), A(10) => 
                           DATA2(10), A(9) => DATA2(9), A(8) => DATA2(8), A(7) 
                           => DATA2(7), A(6) => DATA2(6), A(5) => DATA2(5), 
                           A(4) => DATA2(4), A(3) => DATA2(3), A(2) => DATA2(2)
                           , A(1) => DATA2(1), A(0) => DATA2(0), B(31) => 
                           DATA1(31), B(30) => DATA1(30), B(29) => DATA1(29), 
                           B(28) => DATA1(28), B(27) => DATA1(27), B(26) => 
                           DATA1(26), B(25) => DATA1(25), B(24) => DATA1(24), 
                           B(23) => DATA1(23), B(22) => DATA1(22), B(21) => 
                           DATA1(21), B(20) => DATA1(20), B(19) => DATA1(19), 
                           B(18) => DATA1(18), B(17) => DATA1(17), B(16) => 
                           DATA1(16), B(15) => DATA1(15), B(14) => DATA1(14), 
                           B(13) => DATA1(13), B(12) => DATA1(12), B(11) => 
                           DATA1(11), B(10) => DATA1(10), B(9) => DATA1(9), 
                           B(8) => DATA1(8), B(7) => DATA1(7), B(6) => DATA1(6)
                           , B(5) => DATA1(5), B(4) => DATA1(4), B(3) => 
                           DATA1(3), B(2) => DATA1(2), B(1) => DATA1(1), B(0) 
                           => DATA1(0), TC => n98, LT => n_4441, GT => n_4442, 
                           EQ => n_4443, LE => N2513, GE => N2514, NE => n_4444
                           );
   U3 : OR2_X1 port map( A1 => n1022, A2 => n375, ZN => n2);
   U4 : OR2_X1 port map( A1 => n1032, A2 => DATA2(0), ZN => n3);
   U6 : OR3_X1 port map( A1 => n1034, A2 => n553, A3 => n730, ZN => n4);
   U7 : OR2_X1 port map( A1 => n247, A2 => n1031, ZN => n5);
   U8 : OR2_X1 port map( A1 => n15, A2 => n1027, ZN => n6);
   U9 : NOR2_X2 port map( A1 => n252, A2 => n729, ZN => n62);
   U10 : NAND2_X2 port map( A1 => n219, A2 => n10, ZN => n216);
   U11 : INV_X2 port map( A => n316, ZN => n221);
   U12 : INV_X2 port map( A => n554, ZN => n31);
   U13 : NOR2_X4 port map( A1 => n27, A2 => n28, ZN => n554);
   U14 : INV_X2 port map( A => n2, ZN => n7);
   U15 : INV_X2 port map( A => n4, ZN => n8);
   U16 : INV_X1 port map( A => n218, ZN => n9);
   U17 : INV_X2 port map( A => n9, ZN => n10);
   U18 : INV_X1 port map( A => n227, ZN => n11);
   U19 : INV_X2 port map( A => n11, ZN => n12);
   U20 : NAND2_X4 port map( A1 => n1031, A2 => n1032, ZN => n245);
   U21 : INV_X4 port map( A => n534, ZN => n165);
   U22 : NAND2_X4 port map( A1 => n1026, A2 => n980, ZN => n247);
   U23 : OR2_X1 port map( A1 => n15, A2 => n16, ZN => n139);
   U24 : INV_X4 port map( A => n139, ZN => n13);
   U25 : INV_X1 port map( A => n242, ZN => n14);
   U26 : INV_X4 port map( A => n14, ZN => n15);
   U27 : INV_X4 port map( A => n6, ZN => n16);
   U28 : INV_X4 port map( A => n5, ZN => n17);
   U29 : INV_X4 port map( A => n3, ZN => n18);
   U30 : AND3_X2 port map( A1 => n723, A2 => n726, A3 => n728, ZN => n28);
   U31 : AND3_X2 port map( A1 => n728, A2 => n726, A3 => FUNC(3), ZN => n27);
   U32 : NAND2_X2 port map( A1 => n617, A2 => n970, ZN => n205);
   U33 : OAI21_X2 port map( B1 => n773, B2 => n780, A => n192, ZN => n111);
   U34 : AOI21_X2 port map( B1 => DATA2(4), B2 => n859, A => n1033, ZN => n192)
                           ;
   U35 : NAND3_X2 port map( A1 => n723, A2 => n726, A3 => n727, ZN => n83);
   U36 : NAND2_X2 port map( A1 => n1022, A2 => n1023, ZN => n94);
   U37 : OAI21_X4 port map( B1 => DATA2(0), B2 => n979, A => n971, ZN => n212);
   U38 : NOR2_X4 port map( A1 => n1011, A2 => n1010, ZN => n223);
   U39 : NAND3_X2 port map( A1 => n728, A2 => n723, A3 => FUNC(2), ZN => n553);
   U40 : NAND2_X2 port map( A1 => n1011, A2 => n764, ZN => n375);
   U41 : INV_X2 port map( A => n274, ZN => n228);
   U42 : NAND2_X2 port map( A1 => n228, A2 => n1010, ZN => n231);
   U43 : NOR2_X2 port map( A1 => n922, A2 => n924, ZN => n78);
   U44 : NAND2_X2 port map( A1 => n1026, A2 => n65, ZN => n92);
   U45 : NAND2_X2 port map( A1 => n727, A2 => n726, ZN => n84);
   U46 : AOI21_X4 port map( B1 => DATA2(1), B2 => n1027, A => n1023, ZN => n376
                           );
   U47 : NOR2_X4 port map( A1 => DATA2(5), A2 => DATA2(4), ZN => n219);
   U48 : AOI21_X1 port map( B1 => n19, B2 => n20, A => n553, ZN => 
                           zero_mul_detect);
   U49 : MUX2_X1 port map( A => n21, B => n22, S => signed_notsigned, Z => 
                           overflow);
   U50 : NOR2_X1 port map( A1 => n23, A2 => n24, ZN => n22);
   U51 : MUX2_X1 port map( A => n25, B => n26, S => adder_out_31_port, Z => n23
                           );
   U52 : AOI22_X1 port map( A1 => n27, A2 => DATA2(31), B1 => n28, B2 => n29, 
                           ZN => n26);
   U53 : AOI22_X1 port map( A1 => n27, A2 => n30, B1 => n28, B2 => DATA1(31), 
                           ZN => n25);
   U54 : AND2_X1 port map( A1 => cout, A2 => n31, ZN => n21);
   U55 : AOI21_X1 port map( B1 => n32, B2 => n33, A => n553, ZN => 
                           mul_exeception);
   U56 : NOR4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           n33);
   U57 : OR4_X1 port map( A1 => DATA1(31), A2 => DATA2(16), A3 => DATA2(17), A4
                           => DATA2(18), ZN => n37);
   U58 : OR4_X1 port map( A1 => DATA2(19), A2 => DATA2(20), A3 => DATA2(21), A4
                           => DATA2(22), ZN => n36);
   U59 : OR4_X1 port map( A1 => DATA2(23), A2 => DATA2(24), A3 => DATA2(25), A4
                           => DATA2(26), ZN => n35);
   U60 : OR4_X1 port map( A1 => DATA2(30), A2 => DATA2(31), A3 => DATA2(29), A4
                           => n38, ZN => n34);
   U61 : OR2_X1 port map( A1 => DATA2(28), A2 => DATA2(27), ZN => n38);
   U62 : NOR4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           n32);
   U63 : NAND4_X1 port map( A1 => check_mul_logic, A2 => n43, A3 => n44, A4 => 
                           n45, ZN => n42);
   U64 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           n41);
   U65 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           n40);
   U66 : NAND4_X1 port map( A1 => n54, A2 => n55, A3 => n56, A4 => n57, ZN => 
                           n39);
   U67 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => OUTALU(9));
   U68 : AOI222_X1 port map( A1 => dataout_mul_9_port, A2 => n8, B1 => n60, B2 
                           => n61, C1 => n62, C2 => n63, ZN => n59);
   U69 : OAI221_X1 port map( B1 => n64, B2 => n65, C1 => n66, C2 => n2, A => 
                           n67, ZN => n63);
   U70 : AOI22_X1 port map( A1 => n68, A2 => n69, B1 => n70, B2 => n71, ZN => 
                           n67);
   U71 : INV_X1 port map( A => n72, ZN => n61);
   U72 : AOI222_X1 port map( A1 => n73, A2 => n74, B1 => n75, B2 => n76, C1 => 
                           n77, C2 => n78, ZN => n72);
   U73 : AOI21_X1 port map( B1 => adder_out_9_port, B2 => n31, A => n79, ZN => 
                           n58);
   U74 : MUX2_X1 port map( A => n80, B => n81, S => DATA2(9), Z => n79);
   U75 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => n81);
   U76 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(9), Z => n82);
   U77 : NOR2_X1 port map( A1 => n84, A2 => n86, ZN => n80);
   U78 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => OUTALU(8));
   U79 : AOI222_X1 port map( A1 => dataout_mul_8_port, A2 => n8, B1 => n60, B2 
                           => n89, C1 => n62, C2 => n90, ZN => n88);
   U80 : OAI222_X1 port map( A1 => n91, A2 => n92, B1 => n93, B2 => n65, C1 => 
                           n66, C2 => n94, ZN => n90);
   U81 : OAI221_X1 port map( B1 => n95, B2 => n96, C1 => n97, C2 => n99, A => 
                           n100, ZN => n89);
   U82 : AOI22_X1 port map( A1 => n74, A2 => n75, B1 => n78, B2 => n73, ZN => 
                           n100);
   U83 : INV_X1 port map( A => n101, ZN => n95);
   U84 : AOI21_X1 port map( B1 => adder_out_8_port, B2 => n31, A => n102, ZN =>
                           n87);
   U85 : MUX2_X1 port map( A => n103, B => n104, S => DATA2(8), Z => n102);
   U86 : NAND2_X1 port map( A1 => n105, A2 => n83, ZN => n104);
   U87 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(8), Z => n105);
   U88 : NOR2_X1 port map( A1 => n84, A2 => n106, ZN => n103);
   U89 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => OUTALU(7));
   U90 : AOI221_X1 port map( B1 => dataout_mul_7_port, B2 => n8, C1 => n62, C2 
                           => n109, A => n110, ZN => n108);
   U91 : NOR3_X1 port map( A1 => n111, A2 => n112, A3 => n113, ZN => n110);
   U92 : OAI22_X1 port map( A1 => n66, A2 => n92, B1 => n91, B2 => n65, ZN => 
                           n109);
   U93 : AOI21_X1 port map( B1 => adder_out_7_port, B2 => n31, A => n114, ZN =>
                           n107);
   U94 : MUX2_X1 port map( A => n115, B => n116, S => DATA2(7), Z => n114);
   U95 : NAND2_X1 port map( A1 => n117, A2 => n83, ZN => n116);
   U96 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(7), Z => n117);
   U97 : NOR2_X1 port map( A1 => n84, A2 => n118, ZN => n115);
   U98 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => OUTALU(6));
   U99 : AOI221_X1 port map( B1 => dataout_mul_6_port, B2 => n8, C1 => n60, C2 
                           => n121, A => n122, ZN => n120);
   U100 : NOR3_X1 port map( A1 => n123, A2 => n66, A3 => n65, ZN => n122);
   U101 : OAI22_X1 port map( A1 => n124, A2 => n111, B1 => n112, B2 => n125, ZN
                           => n121);
   U103 : AOI21_X1 port map( B1 => adder_out_6_port, B2 => n31, A => n126, ZN 
                           => n119);
   U104 : MUX2_X1 port map( A => n127, B => n128, S => DATA2(6), Z => n126);
   U105 : NAND2_X1 port map( A1 => n129, A2 => n83, ZN => n128);
   U106 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(6), Z => n129);
   U107 : NOR2_X1 port map( A1 => n84, A2 => n130, ZN => n127);
   U108 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => OUTALU(5));
   U109 : AOI221_X1 port map( B1 => dataout_mul_5_port, B2 => n8, C1 => n62, C2
                           => n133, A => n134, ZN => n132);
   U110 : NOR3_X1 port map( A1 => n135, A2 => n136, A3 => n113, ZN => n134);
   U111 : INV_X1 port map( A => n137, ZN => n133);
   U112 : AOI22_X1 port map( A1 => n138, A2 => n13, B1 => n140, B2 => n16, ZN 
                           => n137);
   U113 : AOI21_X1 port map( B1 => adder_out_5_port, B2 => n31, A => n141, ZN 
                           => n131);
   U114 : MUX2_X1 port map( A => n142, B => n143, S => DATA2(5), Z => n141);
   U115 : NAND2_X1 port map( A1 => n144, A2 => n83, ZN => n143);
   U116 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(5), Z => n144);
   U117 : NOR2_X1 port map( A1 => n84, A2 => n145, ZN => n142);
   U118 : NAND2_X1 port map( A1 => n146, A2 => n147, ZN => OUTALU(4));
   U119 : AOI221_X1 port map( B1 => dataout_mul_4_port, B2 => n8, C1 => n60, C2
                           => n148, A => n149, ZN => n147);
   U120 : AND3_X1 port map( A1 => n62, A2 => n138, A3 => n16, ZN => n149);
   U121 : OAI22_X1 port map( A1 => n136, A2 => n150, B1 => n151, B2 => n135, ZN
                           => n148);
   U122 : AOI21_X1 port map( B1 => adder_out_4_port, B2 => n31, A => n152, ZN 
                           => n146);
   U123 : MUX2_X1 port map( A => n153, B => n154, S => DATA2(4), Z => n152);
   U124 : NAND2_X1 port map( A1 => n155, A2 => n83, ZN => n154);
   U125 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(4), Z => n155);
   U126 : NOR2_X1 port map( A1 => n84, A2 => n156, ZN => n153);
   U127 : NAND2_X1 port map( A1 => n157, A2 => n158, ZN => OUTALU(3));
   U128 : AOI222_X1 port map( A1 => dataout_mul_3_port, A2 => n8, B1 => n62, B2
                           => n159, C1 => n60, C2 => n160, ZN => n158);
   U129 : OAI222_X1 port map( A1 => n151, A2 => n150, B1 => n161, B2 => n135, 
                           C1 => n136, C2 => n162, ZN => n160);
   U130 : INV_X1 port map( A => n163, ZN => n151);
   U131 : OAI221_X1 port map( B1 => n3, B2 => n164, C1 => n165, C2 => n166, A 
                           => n167, ZN => n159);
   U132 : AOI22_X1 port map( A1 => DATA1(0), A2 => n17, B1 => DATA1(1), B2 => 
                           n168, ZN => n167);
   U133 : AOI21_X1 port map( B1 => adder_out_3_port, B2 => n31, A => n169, ZN 
                           => n157);
   U134 : MUX2_X1 port map( A => n170, B => n171, S => DATA2(3), Z => n169);
   U135 : NAND2_X1 port map( A1 => n172, A2 => n83, ZN => n171);
   U136 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(3), Z => n172);
   U137 : NOR2_X1 port map( A1 => n84, A2 => n164, ZN => n170);
   U138 : NAND2_X1 port map( A1 => n173, A2 => n174, ZN => OUTALU(31));
   U139 : AOI221_X1 port map( B1 => DATA2(31), B2 => n175, C1 => n176, C2 => 
                           n60, A => n177, ZN => n174);
   U140 : OAI22_X1 port map( A1 => n24, A2 => n84, B1 => n178, B2 => n123, ZN 
                           => n177);
   U141 : AOI221_X1 port map( B1 => n179, B2 => n180, C1 => n181, C2 => n182, A
                           => n183, ZN => n178);
   U142 : INV_X1 port map( A => n184, ZN => n183);
   U143 : AOI222_X1 port map( A1 => n185, A2 => n186, B1 => n187, B2 => n188, 
                           C1 => n189, C2 => n190, ZN => n184);
   U144 : OAI222_X1 port map( A1 => n191, A2 => n192, B1 => n111, B2 => n193, 
                           C1 => n125, C2 => n194, ZN => n187);
   U145 : AOI221_X1 port map( B1 => n195, B2 => n74, C1 => n196, C2 => n78, A 
                           => n197, ZN => n193);
   U146 : INV_X1 port map( A => n198, ZN => n197);
   U147 : AOI222_X1 port map( A1 => n199, A2 => n200, B1 => n201, B2 => n202, 
                           C1 => n76, C2 => n203, ZN => n198);
   U148 : OAI221_X1 port map( B1 => n204, B2 => n205, C1 => n206, C2 => n207, A
                           => n208, ZN => n203);
   U149 : AOI222_X1 port map( A1 => n209, A2 => n210, B1 => n211, B2 => n212, 
                           C1 => n213, C2 => n214, ZN => n208);
   U150 : OAI222_X1 port map( A1 => n215, A2 => n216, B1 => n217, B2 => n10, C1
                           => n219, C2 => n220, ZN => n211);
   U151 : AOI221_X1 port map( B1 => n221, B2 => n222, C1 => n223, C2 => n224, A
                           => n225, ZN => n217);
   U152 : OAI222_X1 port map( A1 => n226, A2 => n12, B1 => n228, B2 => n229, C1
                           => n230, C2 => n231, ZN => n225);
   U153 : INV_X1 port map( A => n232, ZN => n226);
   U154 : OAI221_X1 port map( B1 => n92, B2 => n233, C1 => n94, C2 => n234, A 
                           => n235, ZN => n232);
   U155 : INV_X1 port map( A => n236, ZN => n235);
   U156 : OAI222_X1 port map( A1 => n237, A2 => n238, B1 => n239, B2 => n65, C1
                           => n240, C2 => n2, ZN => n236);
   U157 : AOI222_X1 port map( A1 => n241, A2 => n15, B1 => n16, B2 => n243, C1 
                           => n13, C2 => n244, ZN => n239);
   U158 : OAI221_X1 port map( B1 => n165, B2 => n57, C1 => n56, C2 => n245, A 
                           => n246, ZN => n243);
   U159 : AOI221_X1 port map( B1 => DATA1(28), B2 => n17, C1 => DATA1(27), C2 
                           => n247, A => n176, ZN => n246);
   U160 : INV_X1 port map( A => n248, ZN => n204);
   U161 : XOR2_X1 port map( A => n30, B => DATA1(31), Z => n24);
   U162 : INV_X1 port map( A => DATA2(31), ZN => n30);
   U163 : NOR2_X1 port map( A1 => n29, A2 => n3, ZN => n176);
   U164 : OAI21_X1 port map( B1 => n29, B2 => n85, A => n83, ZN => n175);
   U165 : AOI221_X1 port map( B1 => adder_out_31_port, B2 => n31, C1 => 
                           dataout_mul_31_port, C2 => n8, A => n249, ZN => n173
                           );
   U166 : NOR4_X1 port map( A1 => DATA2(5), A2 => n250, A3 => n251, A4 => n252,
                           ZN => n249);
   U167 : NAND2_X1 port map( A1 => n253, A2 => n254, ZN => OUTALU(30));
   U168 : AOI222_X1 port map( A1 => dataout_mul_30_port, A2 => n8, B1 => n62, 
                           B2 => n255, C1 => n60, C2 => n256, ZN => n254);
   U169 : OAI22_X1 port map( A1 => n29, A2 => n165, B1 => n3, B2 => n57, ZN => 
                           n256);
   U170 : INV_X1 port map( A => n251, ZN => n255);
   U171 : AOI221_X1 port map( B1 => n182, B2 => n179, C1 => n189, C2 => n181, A
                           => n257, ZN => n251);
   U172 : INV_X1 port map( A => n258, ZN => n257);
   U173 : AOI222_X1 port map( A1 => n190, A2 => n185, B1 => n186, B2 => n259, 
                           C1 => n188, C2 => n180, ZN => n258);
   U174 : OAI222_X1 port map( A1 => n191, A2 => n125, B1 => n194, B2 => n111, 
                           C1 => n192, C2 => n260, ZN => n180);
   U175 : AOI221_X1 port map( B1 => n196, B2 => n74, C1 => n200, C2 => n78, A 
                           => n261, ZN => n194);
   U176 : INV_X1 port map( A => n262, ZN => n261);
   U177 : AOI222_X1 port map( A1 => n199, A2 => n202, B1 => n201, B2 => n263, 
                           C1 => n76, C2 => n195, ZN => n262);
   U178 : OAI221_X1 port map( B1 => n206, B2 => n205, C1 => n264, C2 => n207, A
                           => n265, ZN => n195);
   U179 : AOI222_X1 port map( A1 => n209, A2 => n213, B1 => n266, B2 => n214, 
                           C1 => n248, C2 => n212, ZN => n265);
   U180 : OAI222_X1 port map( A1 => n220, A2 => n216, B1 => n215, B2 => n10, C1
                           => n219, C2 => n267, ZN => n248);
   U181 : AOI221_X1 port map( B1 => n224, B2 => n221, C1 => n268, C2 => n223, A
                           => n269, ZN => n215);
   U182 : INV_X1 port map( A => n270, ZN => n269);
   U183 : AOI222_X1 port map( A1 => n271, A2 => n272, B1 => n273, B2 => n274, 
                           C1 => n11, C2 => n222, ZN => n270);
   U184 : OAI221_X1 port map( B1 => n234, B2 => n92, C1 => n240, C2 => n94, A 
                           => n275, ZN => n222);
   U185 : INV_X1 port map( A => n276, ZN => n275);
   U186 : OAI222_X1 port map( A1 => n2, A2 => n238, B1 => n277, B2 => n237, C1 
                           => n65, C2 => n233, ZN => n276);
   U187 : AOI222_X1 port map( A1 => n241, A2 => n13, B1 => n244, B2 => n16, C1 
                           => n15, C2 => n278, ZN => n233);
   U188 : OAI221_X1 port map( B1 => n56, B2 => n165, C1 => n55, C2 => n245, A 
                           => n279, ZN => n244);
   U189 : AOI222_X1 port map( A1 => DATA1(27), A2 => n17, B1 => DATA1(26), B2 
                           => n247, C1 => DATA1(30), C2 => n18, ZN => n279);
   U190 : INV_X1 port map( A => n230, ZN => n268);
   U191 : INV_X1 port map( A => n280, ZN => n206);
   U192 : AOI21_X1 port map( B1 => adder_out_30_port, B2 => n31, A => n281, ZN 
                           => n253);
   U193 : MUX2_X1 port map( A => n282, B => n283, S => DATA2(30), Z => n281);
   U194 : NAND2_X1 port map( A1 => n284, A2 => n83, ZN => n283);
   U195 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(30), Z => n284);
   U196 : NOR2_X1 port map( A1 => n84, A2 => n57, ZN => n282);
   U197 : NAND2_X1 port map( A1 => n285, A2 => n286, ZN => OUTALU(2));
   U198 : AOI222_X1 port map( A1 => dataout_mul_2_port, A2 => n8, B1 => n62, B2
                           => n287, C1 => n60, C2 => n288, ZN => n286);
   U199 : OAI221_X1 port map( B1 => n289, B2 => n135, C1 => n136, C2 => n290, A
                           => n291, ZN => n288);
   U200 : AOI22_X1 port map( A1 => n179, A2 => n292, B1 => n181, B2 => n163, ZN
                           => n291);
   U201 : INV_X1 port map( A => n293, ZN => n136);
   U202 : OAI222_X1 port map( A1 => n294, A2 => n245, B1 => n165, B2 => n295, 
                           C1 => n3, C2 => n166, ZN => n287);
   U203 : AOI21_X1 port map( B1 => adder_out_2_port, B2 => n31, A => n296, ZN 
                           => n285);
   U204 : MUX2_X1 port map( A => n297, B => n298, S => DATA2(2), Z => n296);
   U205 : NAND2_X1 port map( A1 => n299, A2 => n83, ZN => n298);
   U206 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(2), Z => n299);
   U207 : NOR2_X1 port map( A1 => n84, A2 => n166, ZN => n297);
   U208 : NAND2_X1 port map( A1 => n300, A2 => n301, ZN => OUTALU(29));
   U209 : AOI222_X1 port map( A1 => dataout_mul_29_port, A2 => n8, B1 => n62, 
                           B2 => n302, C1 => n60, C2 => n303, ZN => n301);
   U210 : OAI222_X1 port map( A1 => n29, A2 => n245, B1 => n165, B2 => n57, C1 
                           => n3, C2 => n56, ZN => n303);
   U211 : INV_X1 port map( A => DATA1(30), ZN => n57);
   U212 : INV_X1 port map( A => DATA1(31), ZN => n29);
   U213 : INV_X1 port map( A => n304, ZN => n302);
   U214 : AOI221_X1 port map( B1 => n189, B2 => n179, C1 => n185, C2 => n181, A
                           => n305, ZN => n304);
   U215 : INV_X1 port map( A => n306, ZN => n305);
   U216 : AOI22_X1 port map( A1 => n188, A2 => n182, B1 => n190, B2 => n259, ZN
                           => n306);
   U217 : OAI222_X1 port map( A1 => n260, A2 => n125, B1 => n191, B2 => n111, 
                           C1 => n192, C2 => n307, ZN => n182);
   U218 : AOI221_X1 port map( B1 => n200, B2 => n74, C1 => n202, C2 => n78, A 
                           => n308, ZN => n191);
   U219 : INV_X1 port map( A => n309, ZN => n308);
   U220 : AOI222_X1 port map( A1 => n199, A2 => n263, B1 => n201, B2 => n310, 
                           C1 => n76, C2 => n196, ZN => n309);
   U221 : OAI221_X1 port map( B1 => n264, B2 => n205, C1 => n311, C2 => n207, A
                           => n312, ZN => n196);
   U222 : AOI222_X1 port map( A1 => n209, A2 => n266, B1 => n313, B2 => n214, 
                           C1 => n280, C2 => n212, ZN => n312);
   U223 : OAI222_X1 port map( A1 => n267, A2 => n216, B1 => n220, B2 => n10, C1
                           => n219, C2 => n314, ZN => n280);
   U224 : INV_X1 port map( A => n315, ZN => n220);
   U225 : OAI221_X1 port map( B1 => n230, B2 => n316, C1 => n229, C2 => n317, A
                           => n318, ZN => n315);
   U226 : AOI222_X1 port map( A1 => n271, A2 => n273, B1 => n319, B2 => n274, 
                           C1 => n11, C2 => n224, ZN => n318);
   U227 : OAI221_X1 port map( B1 => n240, B2 => n92, C1 => n238, C2 => n94, A 
                           => n320, ZN => n224);
   U228 : INV_X1 port map( A => n321, ZN => n320);
   U229 : OAI222_X1 port map( A1 => n2, A2 => n277, B1 => n322, B2 => n237, C1 
                           => n65, C2 => n234, ZN => n321);
   U230 : AOI222_X1 port map( A1 => n278, A2 => n13, B1 => n241, B2 => n16, C1 
                           => n15, C2 => n323, ZN => n234);
   U231 : OAI221_X1 port map( B1 => n55, B2 => n165, C1 => n245, C2 => n54, A 
                           => n324, ZN => n241);
   U232 : AOI222_X1 port map( A1 => DATA1(26), A2 => n17, B1 => DATA1(25), B2 
                           => n247, C1 => DATA1(29), C2 => n18, ZN => n324);
   U233 : INV_X1 port map( A => n210, ZN => n264);
   U234 : AOI21_X1 port map( B1 => adder_out_29_port, B2 => n31, A => n325, ZN 
                           => n300);
   U235 : MUX2_X1 port map( A => n326, B => n327, S => DATA2(29), Z => n325);
   U236 : NAND2_X1 port map( A1 => n328, A2 => n83, ZN => n327);
   U237 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(29), Z => n328);
   U238 : NOR2_X1 port map( A1 => n84, A2 => n56, ZN => n326);
   U239 : OAI211_X1 port map( C1 => n329, C2 => n123, A => n330, B => n331, ZN 
                           => OUTALU(28));
   U240 : AOI222_X1 port map( A1 => adder_out_28_port, A2 => n31, B1 => n60, B2
                           => n332, C1 => dataout_mul_28_port, C2 => n8, ZN => 
                           n331);
   U241 : OAI221_X1 port map( B1 => n3, B2 => n55, C1 => n56, C2 => n165, A => 
                           n333, ZN => n332);
   U242 : AOI22_X1 port map( A1 => n17, A2 => DATA1(31), B1 => DATA1(30), B2 =>
                           n168, ZN => n333);
   U243 : INV_X1 port map( A => n245, ZN => n168);
   U244 : AOI22_X1 port map( A1 => DATA1(28), A2 => n334, B1 => DATA2(28), B2 
                           => n335, ZN => n330);
   U245 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(28), Z => n335);
   U246 : OAI21_X1 port map( B1 => DATA2(28), B2 => n84, A => n83, ZN => n334);
   U247 : AOI222_X1 port map( A1 => n181, A2 => n259, B1 => n188, B2 => n189, 
                           C1 => n179, C2 => n185, ZN => n329);
   U248 : OAI222_X1 port map( A1 => n307, A2 => n125, B1 => n260, B2 => n111, 
                           C1 => n192, C2 => n338, ZN => n189);
   U249 : AOI221_X1 port map( B1 => n202, B2 => n74, C1 => n263, C2 => n78, A 
                           => n339, ZN => n260);
   U250 : INV_X1 port map( A => n340, ZN => n339);
   U251 : AOI222_X1 port map( A1 => n199, A2 => n310, B1 => n201, B2 => n341, 
                           C1 => n76, C2 => n200, ZN => n340);
   U252 : OAI221_X1 port map( B1 => n311, B2 => n205, C1 => n342, C2 => n207, A
                           => n343, ZN => n200);
   U253 : AOI222_X1 port map( A1 => n209, A2 => n313, B1 => n344, B2 => n214, 
                           C1 => n210, C2 => n212, ZN => n343);
   U254 : OAI222_X1 port map( A1 => n314, A2 => n216, B1 => n267, B2 => n10, C1
                           => n219, C2 => n345, ZN => n210);
   U255 : AOI221_X1 port map( B1 => n272, B2 => n221, C1 => n273, C2 => n223, A
                           => n346, ZN => n267);
   U256 : OAI222_X1 port map( A1 => n231, A2 => n347, B1 => n348, B2 => n228, 
                           C1 => n12, C2 => n230, ZN => n346);
   U257 : AOI221_X1 port map( B1 => n349, B2 => n68, C1 => n350, C2 => n70, A 
                           => n351, ZN => n230);
   U258 : OAI222_X1 port map( A1 => n2, A2 => n322, B1 => n352, B2 => n237, C1 
                           => n65, C2 => n240, ZN => n351);
   U259 : AOI222_X1 port map( A1 => n323, A2 => n13, B1 => n278, B2 => n16, C1 
                           => n15, C2 => n353, ZN => n240);
   U260 : OAI221_X1 port map( B1 => n165, B2 => n54, C1 => n53, C2 => n245, A 
                           => n354, ZN => n278);
   U261 : AOI222_X1 port map( A1 => n17, A2 => DATA1(25), B1 => DATA1(24), B2 
                           => n247, C1 => DATA1(28), C2 => n18, ZN => n354);
   U262 : INV_X1 port map( A => n213, ZN => n311);
   U263 : OAI211_X1 port map( C1 => n355, C2 => n123, A => n356, B => n357, ZN 
                           => OUTALU(27));
   U264 : AOI221_X1 port map( B1 => adder_out_27_port, B2 => n31, C1 => 
                           dataout_mul_27_port, C2 => n8, A => n358, ZN => n357
                           );
   U265 : AND3_X1 port map( A1 => n60, A2 => n359, A3 => n16, ZN => n358);
   U266 : AOI22_X1 port map( A1 => DATA1(27), A2 => n360, B1 => DATA2(27), B2 
                           => n361, ZN => n356);
   U267 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(27), Z => n361);
   U268 : OAI21_X1 port map( B1 => DATA2(27), B2 => n84, A => n83, ZN => n360);
   U269 : AOI22_X1 port map( A1 => n188, A2 => n185, B1 => n179, B2 => n259, ZN
                           => n355);
   U270 : OAI222_X1 port map( A1 => n338, A2 => n125, B1 => n307, B2 => n111, 
                           C1 => n192, C2 => n362, ZN => n185);
   U271 : AOI221_X1 port map( B1 => n263, B2 => n74, C1 => n310, C2 => n78, A 
                           => n363, ZN => n307);
   U272 : INV_X1 port map( A => n364, ZN => n363);
   U273 : AOI222_X1 port map( A1 => n199, A2 => n341, B1 => n201, B2 => n365, 
                           C1 => n76, C2 => n202, ZN => n364);
   U274 : OAI221_X1 port map( B1 => n342, B2 => n205, C1 => n366, C2 => n207, A
                           => n367, ZN => n202);
   U275 : AOI222_X1 port map( A1 => n209, A2 => n344, B1 => n368, B2 => n214, 
                           C1 => n213, C2 => n212, ZN => n367);
   U276 : OAI222_X1 port map( A1 => n345, A2 => n216, B1 => n314, B2 => n10, C1
                           => n219, C2 => n369, ZN => n213);
   U277 : AOI221_X1 port map( B1 => n273, B2 => n221, C1 => n319, C2 => n223, A
                           => n370, ZN => n314);
   U278 : OAI222_X1 port map( A1 => n231, A2 => n348, B1 => n371, B2 => n228, 
                           C1 => n12, C2 => n229, ZN => n370);
   U279 : INV_X1 port map( A => n272, ZN => n229);
   U280 : OAI221_X1 port map( B1 => n277, B2 => n92, C1 => n322, C2 => n94, A 
                           => n372, ZN => n272);
   U281 : AOI222_X1 port map( A1 => n7, A2 => n373, B1 => n374, B2 => n375, C1 
                           => n376, C2 => n349, ZN => n372);
   U282 : INV_X1 port map( A => n238, ZN => n349);
   U283 : AOI222_X1 port map( A1 => n353, A2 => n13, B1 => n323, B2 => n16, C1 
                           => n15, C2 => n377, ZN => n238);
   U284 : OAI221_X1 port map( B1 => n165, B2 => n53, C1 => n52, C2 => n245, A 
                           => n378, ZN => n323);
   U285 : AOI222_X1 port map( A1 => DATA1(24), A2 => n17, B1 => DATA1(23), B2 
                           => n247, C1 => DATA1(27), C2 => n18, ZN => n378);
   U286 : INV_X1 port map( A => n266, ZN => n342);
   U287 : NAND3_X1 port map( A1 => n379, A2 => n380, A3 => n381, ZN => 
                           OUTALU(26));
   U288 : AOI222_X1 port map( A1 => adder_out_26_port, A2 => n31, B1 => n60, B2
                           => n382, C1 => dataout_mul_26_port, C2 => n8, ZN => 
                           n381);
   U289 : INV_X1 port map( A => n383, ZN => n382);
   U290 : AOI22_X1 port map( A1 => n384, A2 => n16, B1 => n359, B2 => n13, ZN 
                           => n383);
   U291 : NAND3_X1 port map( A1 => n62, A2 => n259, A3 => n188, ZN => n380);
   U292 : OAI222_X1 port map( A1 => n362, A2 => n125, B1 => n338, B2 => n111, 
                           C1 => n192, C2 => n385, ZN => n259);
   U293 : AOI221_X1 port map( B1 => n310, B2 => n74, C1 => n341, C2 => n78, A 
                           => n386, ZN => n338);
   U294 : INV_X1 port map( A => n387, ZN => n386);
   U295 : AOI222_X1 port map( A1 => n199, A2 => n365, B1 => n201, B2 => n388, 
                           C1 => n76, C2 => n263, ZN => n387);
   U296 : OAI221_X1 port map( B1 => n366, B2 => n205, C1 => n389, C2 => n207, A
                           => n390, ZN => n263);
   U297 : AOI222_X1 port map( A1 => n209, A2 => n368, B1 => n391, B2 => n214, 
                           C1 => n266, C2 => n212, ZN => n390);
   U298 : OAI222_X1 port map( A1 => n369, A2 => n216, B1 => n345, B2 => n10, C1
                           => n219, C2 => n392, ZN => n266);
   U299 : AOI221_X1 port map( B1 => n319, B2 => n221, C1 => n393, C2 => n223, A
                           => n394, ZN => n345);
   U300 : INV_X1 port map( A => n395, ZN => n394);
   U301 : AOI222_X1 port map( A1 => n271, A2 => n396, B1 => n397, B2 => n274, 
                           C1 => n11, C2 => n273, ZN => n395);
   U302 : OAI221_X1 port map( B1 => n322, B2 => n92, C1 => n352, C2 => n94, A 
                           => n398, ZN => n273);
   U303 : AOI222_X1 port map( A1 => n7, A2 => n374, B1 => n399, B2 => n375, C1 
                           => n376, C2 => n350, ZN => n398);
   U304 : INV_X1 port map( A => n277, ZN => n350);
   U305 : AOI222_X1 port map( A1 => n377, A2 => n13, B1 => n353, B2 => n16, C1 
                           => n15, C2 => n400, ZN => n277);
   U306 : OAI221_X1 port map( B1 => n52, B2 => n165, C1 => n245, C2 => n51, A 
                           => n401, ZN => n353);
   U307 : AOI222_X1 port map( A1 => DATA1(23), A2 => n17, B1 => DATA1(22), B2 
                           => n247, C1 => DATA1(26), C2 => n18, ZN => n401);
   U308 : INV_X1 port map( A => n402, ZN => n399);
   U309 : INV_X1 port map( A => n347, ZN => n319);
   U310 : INV_X1 port map( A => n313, ZN => n366);
   U311 : AOI22_X1 port map( A1 => DATA1(26), A2 => n403, B1 => DATA2(26), B2 
                           => n404, ZN => n379);
   U312 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(26), Z => n404);
   U313 : OAI21_X1 port map( B1 => DATA2(26), B2 => n84, A => n83, ZN => n403);
   U314 : OAI211_X1 port map( C1 => n405, C2 => n123, A => n406, B => n407, ZN 
                           => OUTALU(25));
   U315 : AOI221_X1 port map( B1 => adder_out_25_port, B2 => n31, C1 => 
                           dataout_mul_25_port, C2 => n8, A => n408, ZN => n407
                           );
   U316 : NOR3_X1 port map( A1 => n113, A2 => n409, A3 => n65, ZN => n408);
   U317 : AOI22_X1 port map( A1 => DATA1(25), A2 => n410, B1 => DATA2(25), B2 
                           => n411, ZN => n406);
   U318 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(25), Z => n411);
   U319 : OAI21_X1 port map( B1 => DATA2(25), B2 => n84, A => n83, ZN => n410);
   U320 : INV_X1 port map( A => n412, ZN => n405);
   U321 : OAI22_X1 port map( A1 => n111, A2 => n362, B1 => n125, B2 => n385, ZN
                           => n412);
   U322 : AOI221_X1 port map( B1 => n341, B2 => n74, C1 => n365, C2 => n78, A 
                           => n413, ZN => n362);
   U323 : INV_X1 port map( A => n414, ZN => n413);
   U324 : AOI222_X1 port map( A1 => n199, A2 => n388, B1 => n201, B2 => n415, 
                           C1 => n76, C2 => n310, ZN => n414);
   U325 : OAI221_X1 port map( B1 => n389, B2 => n205, C1 => n416, C2 => n207, A
                           => n417, ZN => n310);
   U326 : AOI222_X1 port map( A1 => n209, A2 => n391, B1 => n418, B2 => n214, 
                           C1 => n313, C2 => n212, ZN => n417);
   U327 : OAI222_X1 port map( A1 => n392, A2 => n216, B1 => n369, B2 => n10, C1
                           => n219, C2 => n419, ZN => n313);
   U328 : AOI221_X1 port map( B1 => n393, B2 => n221, C1 => n396, C2 => n223, A
                           => n420, ZN => n369);
   U329 : OAI222_X1 port map( A1 => n231, A2 => n421, B1 => n422, B2 => n228, 
                           C1 => n12, C2 => n347, ZN => n420);
   U330 : AOI221_X1 port map( B1 => n373, B2 => n68, C1 => n374, C2 => n70, A 
                           => n423, ZN => n347);
   U331 : OAI222_X1 port map( A1 => n2, A2 => n402, B1 => n424, B2 => n237, C1 
                           => n65, C2 => n322, ZN => n423);
   U332 : AOI222_X1 port map( A1 => n400, A2 => n13, B1 => n377, B2 => n16, C1 
                           => n15, C2 => n425, ZN => n322);
   U333 : OAI221_X1 port map( B1 => n165, B2 => n51, C1 => n245, C2 => n50, A 
                           => n426, ZN => n377);
   U334 : AOI222_X1 port map( A1 => DATA1(22), A2 => n17, B1 => DATA1(21), B2 
                           => n247, C1 => DATA1(25), C2 => n18, ZN => n426);
   U335 : INV_X1 port map( A => n344, ZN => n389);
   U336 : NAND3_X1 port map( A1 => n427, A2 => n428, A3 => n429, ZN => 
                           OUTALU(24));
   U337 : AOI222_X1 port map( A1 => adder_out_24_port, A2 => n31, B1 => n60, B2
                           => n430, C1 => dataout_mul_24_port, C2 => n8, ZN => 
                           n429);
   U338 : OAI22_X1 port map( A1 => n409, A2 => n92, B1 => n431, B2 => n65, ZN 
                           => n430);
   U339 : OR3_X1 port map( A1 => n123, A2 => n385, A3 => n111, ZN => n428);
   U340 : AOI221_X1 port map( B1 => n365, B2 => n74, C1 => n388, C2 => n78, A 
                           => n432, ZN => n385);
   U341 : INV_X1 port map( A => n433, ZN => n432);
   U342 : AOI222_X1 port map( A1 => n199, A2 => n415, B1 => n201, B2 => n434, 
                           C1 => n76, C2 => n341, ZN => n433);
   U343 : OAI221_X1 port map( B1 => n416, B2 => n205, C1 => n435, C2 => n207, A
                           => n436, ZN => n341);
   U344 : AOI222_X1 port map( A1 => n209, A2 => n418, B1 => n437, B2 => n214, 
                           C1 => n344, C2 => n212, ZN => n436);
   U345 : OAI222_X1 port map( A1 => n419, A2 => n216, B1 => n392, B2 => n10, C1
                           => n219, C2 => n438, ZN => n344);
   U346 : AOI221_X1 port map( B1 => n396, B2 => n221, C1 => n397, C2 => n223, A
                           => n439, ZN => n392);
   U347 : OAI222_X1 port map( A1 => n231, A2 => n422, B1 => n440, B2 => n228, 
                           C1 => n12, C2 => n348, ZN => n439);
   U348 : INV_X1 port map( A => n393, ZN => n348);
   U349 : OAI221_X1 port map( B1 => n441, B2 => n92, C1 => n402, C2 => n94, A 
                           => n442, ZN => n393);
   U350 : AOI222_X1 port map( A1 => n7, A2 => n443, B1 => n444, B2 => n375, C1 
                           => n376, C2 => n373, ZN => n442);
   U351 : INV_X1 port map( A => n352, ZN => n373);
   U352 : AOI222_X1 port map( A1 => n425, A2 => n13, B1 => n400, B2 => n16, C1 
                           => n15, C2 => n445, ZN => n352);
   U353 : OAI221_X1 port map( B1 => n165, B2 => n50, C1 => n245, C2 => n49, A 
                           => n446, ZN => n400);
   U354 : AOI222_X1 port map( A1 => DATA1(21), A2 => n17, B1 => DATA1(20), B2 
                           => n247, C1 => DATA1(24), C2 => n18, ZN => n446);
   U355 : INV_X1 port map( A => n368, ZN => n416);
   U356 : AOI22_X1 port map( A1 => DATA1(24), A2 => n447, B1 => DATA2(24), B2 
                           => n448, ZN => n427);
   U357 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(24), Z => n448);
   U358 : OAI21_X1 port map( B1 => DATA2(24), B2 => n84, A => n83, ZN => n447);
   U359 : OAI211_X1 port map( C1 => n449, C2 => n123, A => n450, B => n451, ZN 
                           => OUTALU(23));
   U360 : AOI222_X1 port map( A1 => adder_out_23_port, A2 => n31, B1 => n60, B2
                           => n452, C1 => dataout_mul_23_port, C2 => n8, ZN => 
                           n451);
   U361 : OAI222_X1 port map( A1 => n431, A2 => n92, B1 => n453, B2 => n65, C1 
                           => n409, C2 => n94, ZN => n452);
   U362 : AOI22_X1 port map( A1 => DATA1(23), A2 => n454, B1 => DATA2(23), B2 
                           => n455, ZN => n450);
   U363 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(23), Z => n455);
   U364 : OAI21_X1 port map( B1 => DATA2(23), B2 => n84, A => n83, ZN => n454);
   U365 : AOI221_X1 port map( B1 => n74, B2 => n388, C1 => n78, C2 => n415, A 
                           => n456, ZN => n449);
   U366 : INV_X1 port map( A => n457, ZN => n456);
   U367 : AOI22_X1 port map( A1 => n434, A2 => n199, B1 => n365, B2 => n76, ZN 
                           => n457);
   U368 : OAI221_X1 port map( B1 => n435, B2 => n205, C1 => n458, C2 => n207, A
                           => n459, ZN => n365);
   U369 : AOI222_X1 port map( A1 => n209, A2 => n437, B1 => n460, B2 => n214, 
                           C1 => n368, C2 => n212, ZN => n459);
   U370 : OAI222_X1 port map( A1 => n438, A2 => n216, B1 => n419, B2 => n10, C1
                           => n219, C2 => n461, ZN => n368);
   U371 : AOI221_X1 port map( B1 => n397, B2 => n221, C1 => n462, C2 => n223, A
                           => n463, ZN => n419);
   U372 : OAI222_X1 port map( A1 => n231, A2 => n440, B1 => n464, B2 => n228, 
                           C1 => n12, C2 => n371, ZN => n463);
   U373 : INV_X1 port map( A => n396, ZN => n371);
   U374 : OAI221_X1 port map( B1 => n402, B2 => n92, C1 => n424, C2 => n94, A 
                           => n465, ZN => n396);
   U375 : AOI222_X1 port map( A1 => n7, A2 => n444, B1 => n466, B2 => n375, C1 
                           => n376, C2 => n374, ZN => n465);
   U376 : INV_X1 port map( A => n441, ZN => n374);
   U377 : AOI222_X1 port map( A1 => n445, A2 => n13, B1 => n425, B2 => n16, C1 
                           => n15, C2 => n467, ZN => n441);
   U378 : OAI221_X1 port map( B1 => n165, B2 => n49, C1 => n245, C2 => n48, A 
                           => n468, ZN => n425);
   U379 : AOI222_X1 port map( A1 => DATA1(20), A2 => n17, B1 => DATA1(19), B2 
                           => n247, C1 => DATA1(23), C2 => n18, ZN => n468);
   U380 : INV_X1 port map( A => n421, ZN => n397);
   U381 : INV_X1 port map( A => n391, ZN => n435);
   U382 : OAI211_X1 port map( C1 => n469, C2 => n123, A => n470, B => n471, ZN 
                           => OUTALU(22));
   U383 : AOI222_X1 port map( A1 => adder_out_22_port, A2 => n31, B1 => n60, B2
                           => n472, C1 => dataout_mul_22_port, C2 => n8, ZN => 
                           n471);
   U384 : OAI221_X1 port map( B1 => n453, B2 => n92, C1 => n431, C2 => n94, A 
                           => n473, ZN => n472);
   U385 : AOI22_X1 port map( A1 => n376, A2 => n474, B1 => n7, B2 => n475, ZN 
                           => n473);
   U386 : INV_X1 port map( A => n409, ZN => n475);
   U387 : AOI22_X1 port map( A1 => DATA1(22), A2 => n476, B1 => DATA2(22), B2 
                           => n477, ZN => n470);
   U388 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(22), Z => n477);
   U389 : OAI21_X1 port map( B1 => DATA2(22), B2 => n84, A => n83, ZN => n476);
   U390 : AOI222_X1 port map( A1 => n78, A2 => n434, B1 => n76, B2 => n388, C1 
                           => n74, C2 => n415, ZN => n469);
   U391 : OAI221_X1 port map( B1 => n458, B2 => n205, C1 => n478, C2 => n207, A
                           => n479, ZN => n388);
   U392 : AOI222_X1 port map( A1 => n209, A2 => n460, B1 => n480, B2 => n214, 
                           C1 => n391, C2 => n212, ZN => n479);
   U393 : OAI222_X1 port map( A1 => n461, A2 => n216, B1 => n438, B2 => n10, C1
                           => n219, C2 => n481, ZN => n391);
   U394 : AOI221_X1 port map( B1 => n462, B2 => n221, C1 => n482, C2 => n223, A
                           => n483, ZN => n438);
   U395 : OAI222_X1 port map( A1 => n231, A2 => n464, B1 => n484, B2 => n228, 
                           C1 => n12, C2 => n421, ZN => n483);
   U396 : AOI221_X1 port map( B1 => n443, B2 => n68, C1 => n444, C2 => n70, A 
                           => n485, ZN => n421);
   U397 : OAI222_X1 port map( A1 => n2, A2 => n486, B1 => n487, B2 => n237, C1 
                           => n65, C2 => n402, ZN => n485);
   U398 : AOI222_X1 port map( A1 => n467, A2 => n13, B1 => n445, B2 => n16, C1 
                           => n15, C2 => n488, ZN => n402);
   U399 : OAI221_X1 port map( B1 => n165, B2 => n48, C1 => n245, C2 => n47, A 
                           => n489, ZN => n445);
   U400 : AOI222_X1 port map( A1 => DATA1(19), A2 => n17, B1 => DATA1(18), B2 
                           => n247, C1 => DATA1(22), C2 => n18, ZN => n489);
   U401 : INV_X1 port map( A => n418, ZN => n458);
   U402 : OAI211_X1 port map( C1 => n490, C2 => n123, A => n491, B => n492, ZN 
                           => OUTALU(21));
   U403 : AOI221_X1 port map( B1 => adder_out_21_port, B2 => n31, C1 => 
                           dataout_mul_21_port, C2 => n8, A => n493, ZN => n492
                           );
   U404 : NOR3_X1 port map( A1 => n113, A2 => n494, A3 => n12, ZN => n493);
   U405 : AOI22_X1 port map( A1 => DATA1(21), A2 => n495, B1 => DATA2(21), B2 
                           => n496, ZN => n491);
   U406 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(21), Z => n496);
   U407 : OAI21_X1 port map( B1 => DATA2(21), B2 => n84, A => n83, ZN => n495);
   U408 : AOI22_X1 port map( A1 => n76, A2 => n415, B1 => n74, B2 => n434, ZN 
                           => n490);
   U409 : OAI221_X1 port map( B1 => n478, B2 => n205, C1 => n497, C2 => n207, A
                           => n498, ZN => n415);
   U410 : AOI222_X1 port map( A1 => n209, A2 => n480, B1 => n499, B2 => n214, 
                           C1 => n418, C2 => n212, ZN => n498);
   U411 : OAI222_X1 port map( A1 => n481, A2 => n216, B1 => n461, B2 => n10, C1
                           => n219, C2 => n500, ZN => n418);
   U412 : AOI221_X1 port map( B1 => n482, B2 => n221, C1 => n501, C2 => n223, A
                           => n502, ZN => n461);
   U413 : OAI222_X1 port map( A1 => n231, A2 => n484, B1 => n503, B2 => n228, 
                           C1 => n12, C2 => n422, ZN => n502);
   U414 : INV_X1 port map( A => n462, ZN => n422);
   U415 : OAI221_X1 port map( B1 => n504, B2 => n92, C1 => n486, C2 => n94, A 
                           => n505, ZN => n462);
   U416 : AOI222_X1 port map( A1 => n7, A2 => n506, B1 => n507, B2 => n375, C1 
                           => n376, C2 => n443, ZN => n505);
   U417 : INV_X1 port map( A => n424, ZN => n443);
   U418 : AOI222_X1 port map( A1 => n488, A2 => n13, B1 => n467, B2 => n16, C1 
                           => n15, C2 => n508, ZN => n424);
   U419 : OAI221_X1 port map( B1 => n165, B2 => n47, C1 => n245, C2 => n46, A 
                           => n509, ZN => n467);
   U420 : AOI222_X1 port map( A1 => DATA1(18), A2 => n17, B1 => DATA1(17), B2 
                           => n247, C1 => DATA1(21), C2 => n18, ZN => n509);
   U421 : INV_X1 port map( A => n437, ZN => n478);
   U422 : NAND3_X1 port map( A1 => n510, A2 => n511, A3 => n512, ZN => 
                           OUTALU(20));
   U423 : AOI222_X1 port map( A1 => adder_out_20_port, A2 => n31, B1 => n60, B2
                           => n513, C1 => dataout_mul_20_port, C2 => n8, ZN => 
                           n512);
   U424 : OAI22_X1 port map( A1 => n494, A2 => n316, B1 => n514, B2 => n12, ZN 
                           => n513);
   U425 : NAND3_X1 port map( A1 => n76, A2 => n434, A3 => n62, ZN => n511);
   U426 : OAI221_X1 port map( B1 => n497, B2 => n205, C1 => n515, C2 => n207, A
                           => n516, ZN => n434);
   U427 : AOI222_X1 port map( A1 => n209, A2 => n499, B1 => n517, B2 => n214, 
                           C1 => n437, C2 => n212, ZN => n516);
   U428 : OAI222_X1 port map( A1 => n500, A2 => n216, B1 => n481, B2 => n10, C1
                           => n219, C2 => n518, ZN => n437);
   U429 : AOI221_X1 port map( B1 => n501, B2 => n221, C1 => n519, C2 => n223, A
                           => n520, ZN => n481);
   U430 : OAI222_X1 port map( A1 => n231, A2 => n503, B1 => n521, B2 => n228, 
                           C1 => n12, C2 => n440, ZN => n520);
   U431 : INV_X1 port map( A => n482, ZN => n440);
   U432 : OAI221_X1 port map( B1 => n486, B2 => n92, C1 => n487, C2 => n94, A 
                           => n522, ZN => n482);
   U433 : AOI222_X1 port map( A1 => n7, A2 => n507, B1 => n523, B2 => n375, C1 
                           => n376, C2 => n444, ZN => n522);
   U434 : INV_X1 port map( A => n504, ZN => n444);
   U435 : AOI222_X1 port map( A1 => n508, A2 => n13, B1 => n488, B2 => n16, C1 
                           => n15, C2 => n524, ZN => n504);
   U436 : OAI221_X1 port map( B1 => n165, B2 => n46, C1 => n245, C2 => n45, A 
                           => n525, ZN => n488);
   U437 : AOI222_X1 port map( A1 => DATA1(17), A2 => n17, B1 => DATA1(16), B2 
                           => n247, C1 => DATA1(20), C2 => n18, ZN => n525);
   U438 : INV_X1 port map( A => n460, ZN => n497);
   U439 : AOI22_X1 port map( A1 => DATA1(20), A2 => n526, B1 => DATA2(20), B2 
                           => n527, ZN => n510);
   U440 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(20), Z => n527);
   U441 : OAI21_X1 port map( B1 => DATA2(20), B2 => n84, A => n83, ZN => n526);
   U442 : OAI211_X1 port map( C1 => n528, C2 => n123, A => n529, B => n530, ZN 
                           => OUTALU(1));
   U443 : AOI222_X1 port map( A1 => adder_out_1_port, A2 => n31, B1 => n60, B2 
                           => n531, C1 => dataout_mul_1_port, C2 => n8, ZN => 
                           n530);
   U444 : AOI22_X1 port map( A1 => DATA1(1), A2 => n532, B1 => DATA2(1), B2 => 
                           n533, ZN => n529);
   U445 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(1), Z => n533);
   U446 : OAI21_X1 port map( B1 => DATA2(1), B2 => n84, A => n83, ZN => n532);
   U447 : AOI22_X1 port map( A1 => DATA1(0), A2 => n534, B1 => DATA1(1), B2 => 
                           n18, ZN => n528);
   U448 : OAI211_X1 port map( C1 => n535, C2 => n123, A => n536, B => n537, ZN 
                           => OUTALU(19));
   U449 : AOI222_X1 port map( A1 => adder_out_19_port, A2 => n31, B1 => n60, B2
                           => n538, C1 => dataout_mul_19_port, C2 => n8, ZN => 
                           n537);
   U450 : OAI222_X1 port map( A1 => n514, A2 => n316, B1 => n539, B2 => n12, C1
                           => n494, C2 => n317, ZN => n538);
   U451 : AOI22_X1 port map( A1 => DATA1(19), A2 => n540, B1 => DATA2(19), B2 
                           => n541, ZN => n536);
   U452 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(19), Z => n541);
   U453 : OAI21_X1 port map( B1 => DATA2(19), B2 => n84, A => n83, ZN => n540);
   U454 : AOI221_X1 port map( B1 => n460, B2 => n212, C1 => n209, C2 => n517, A
                           => n542, ZN => n535);
   U455 : OAI22_X1 port map( A1 => n543, A2 => n207, B1 => n515, B2 => n205, ZN
                           => n542);
   U456 : INV_X1 port map( A => n480, ZN => n515);
   U457 : INV_X1 port map( A => n499, ZN => n543);
   U458 : OAI222_X1 port map( A1 => n518, A2 => n216, B1 => n500, B2 => n10, C1
                           => n219, C2 => n544, ZN => n460);
   U459 : AOI221_X1 port map( B1 => n519, B2 => n221, C1 => n545, C2 => n223, A
                           => n546, ZN => n500);
   U460 : OAI222_X1 port map( A1 => n231, A2 => n521, B1 => n547, B2 => n228, 
                           C1 => n12, C2 => n464, ZN => n546);
   U461 : INV_X1 port map( A => n501, ZN => n464);
   U462 : OAI221_X1 port map( B1 => n487, B2 => n92, C1 => n548, C2 => n94, A 
                           => n549, ZN => n501);
   U463 : AOI222_X1 port map( A1 => n7, A2 => n523, B1 => n550, B2 => n375, C1 
                           => n376, C2 => n466, ZN => n549);
   U464 : INV_X1 port map( A => n486, ZN => n466);
   U465 : AOI222_X1 port map( A1 => n524, A2 => n13, B1 => n508, B2 => n16, C1 
                           => n15, C2 => n551, ZN => n486);
   U466 : OAI221_X1 port map( B1 => n165, B2 => n45, C1 => n245, C2 => n44, A 
                           => n552, ZN => n508);
   U467 : AOI222_X1 port map( A1 => DATA1(16), A2 => n17, B1 => DATA1(15), B2 
                           => n247, C1 => DATA1(19), C2 => n18, ZN => n552);
   U468 : OAI211_X1 port map( C1 => n555, C2 => n123, A => n556, B => n557, ZN 
                           => OUTALU(18));
   U469 : AOI222_X1 port map( A1 => adder_out_18_port, A2 => n31, B1 => n60, B2
                           => n558, C1 => dataout_mul_18_port, C2 => n8, ZN => 
                           n557);
   U470 : OAI221_X1 port map( B1 => n559, B2 => n12, C1 => n494, C2 => n231, A 
                           => n560, ZN => n558);
   U471 : INV_X1 port map( A => n561, ZN => n560);
   U472 : OAI22_X1 port map( A1 => n316, A2 => n539, B1 => n317, B2 => n514, ZN
                           => n561);
   U473 : AOI22_X1 port map( A1 => DATA1(18), A2 => n562, B1 => DATA2(18), B2 
                           => n563, ZN => n556);
   U474 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(18), Z => n563);
   U475 : OAI21_X1 port map( B1 => DATA2(18), B2 => n84, A => n83, ZN => n562);
   U476 : AOI222_X1 port map( A1 => n564, A2 => n517, B1 => n480, B2 => n212, 
                           C1 => n565, C2 => n499, ZN => n555);
   U477 : OAI222_X1 port map( A1 => n544, A2 => n216, B1 => n518, B2 => n10, C1
                           => n219, C2 => n566, ZN => n480);
   U478 : AOI221_X1 port map( B1 => n545, B2 => n221, C1 => n567, C2 => n223, A
                           => n568, ZN => n518);
   U479 : OAI222_X1 port map( A1 => n231, A2 => n547, B1 => n569, B2 => n228, 
                           C1 => n12, C2 => n484, ZN => n568);
   U480 : INV_X1 port map( A => n519, ZN => n484);
   U481 : OAI221_X1 port map( B1 => n548, B2 => n92, C1 => n570, C2 => n94, A 
                           => n571, ZN => n519);
   U482 : AOI222_X1 port map( A1 => n7, A2 => n550, B1 => n572, B2 => n375, C1 
                           => n376, C2 => n506, ZN => n571);
   U483 : INV_X1 port map( A => n487, ZN => n506);
   U484 : AOI222_X1 port map( A1 => n551, A2 => n13, B1 => n524, B2 => n16, C1 
                           => n15, C2 => n573, ZN => n487);
   U485 : OAI221_X1 port map( B1 => n165, B2 => n44, C1 => n245, C2 => n43, A 
                           => n574, ZN => n524);
   U486 : AOI222_X1 port map( A1 => DATA1(15), A2 => n17, B1 => DATA1(14), B2 
                           => n247, C1 => DATA1(18), C2 => n18, ZN => n574);
   U487 : NAND2_X1 port map( A1 => n575, A2 => n576, ZN => OUTALU(17));
   U488 : AOI221_X1 port map( B1 => dataout_mul_17_port, B2 => n8, C1 => n62, 
                           C2 => n577, A => n578, ZN => n576);
   U489 : NOR3_X1 port map( A1 => n113, A2 => n579, A3 => n10, ZN => n578);
   U490 : INV_X1 port map( A => n580, ZN => n577);
   U491 : AOI22_X1 port map( A1 => n517, A2 => n565, B1 => n212, B2 => n499, ZN
                           => n580);
   U492 : OAI222_X1 port map( A1 => n566, A2 => n216, B1 => n544, B2 => n10, C1
                           => n219, C2 => n581, ZN => n499);
   U493 : AOI221_X1 port map( B1 => n567, B2 => n221, C1 => n582, C2 => n223, A
                           => n583, ZN => n544);
   U494 : OAI222_X1 port map( A1 => n231, A2 => n569, B1 => n584, B2 => n228, 
                           C1 => n12, C2 => n503, ZN => n583);
   U495 : INV_X1 port map( A => n545, ZN => n503);
   U496 : OAI221_X1 port map( B1 => n570, B2 => n92, C1 => n585, C2 => n94, A 
                           => n586, ZN => n545);
   U497 : AOI222_X1 port map( A1 => n7, A2 => n572, B1 => n587, B2 => n375, C1 
                           => n376, C2 => n507, ZN => n586);
   U498 : INV_X1 port map( A => n548, ZN => n507);
   U499 : AOI222_X1 port map( A1 => n573, A2 => n13, B1 => n551, B2 => n16, C1 
                           => n15, C2 => n588, ZN => n548);
   U500 : OAI221_X1 port map( B1 => n165, B2 => n43, C1 => n245, C2 => n589, A 
                           => n590, ZN => n551);
   U501 : AOI222_X1 port map( A1 => DATA1(14), A2 => n17, B1 => DATA1(13), B2 
                           => n247, C1 => DATA1(17), C2 => n18, ZN => n590);
   U502 : AOI21_X1 port map( B1 => adder_out_17_port, B2 => n31, A => n591, ZN 
                           => n575);
   U503 : MUX2_X1 port map( A => n592, B => n593, S => DATA2(17), Z => n591);
   U504 : NAND2_X1 port map( A1 => n594, A2 => n83, ZN => n593);
   U505 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(17), Z => n594);
   U506 : NOR2_X1 port map( A1 => n84, A2 => n44, ZN => n592);
   U507 : NAND3_X1 port map( A1 => n595, A2 => n596, A3 => n597, ZN => 
                           OUTALU(16));
   U508 : AOI222_X1 port map( A1 => adder_out_16_port, A2 => n31, B1 => n60, B2
                           => n598, C1 => dataout_mul_16_port, C2 => n8, ZN => 
                           n597);
   U509 : OAI22_X1 port map( A1 => n579, A2 => n216, B1 => n599, B2 => n10, ZN 
                           => n598);
   U510 : NAND3_X1 port map( A1 => n517, A2 => n212, A3 => n62, ZN => n596);
   U511 : OAI222_X1 port map( A1 => n581, A2 => n216, B1 => n566, B2 => n10, C1
                           => n219, C2 => n600, ZN => n517);
   U512 : AOI221_X1 port map( B1 => n582, B2 => n221, C1 => n601, C2 => n223, A
                           => n602, ZN => n566);
   U513 : OAI222_X1 port map( A1 => n231, A2 => n584, B1 => n603, B2 => n228, 
                           C1 => n12, C2 => n521, ZN => n602);
   U514 : INV_X1 port map( A => n567, ZN => n521);
   U515 : OAI221_X1 port map( B1 => n585, B2 => n92, C1 => n604, C2 => n94, A 
                           => n605, ZN => n567);
   U516 : AOI222_X1 port map( A1 => n7, A2 => n587, B1 => n606, B2 => n375, C1 
                           => n376, C2 => n523, ZN => n605);
   U517 : INV_X1 port map( A => n570, ZN => n523);
   U518 : AOI222_X1 port map( A1 => n588, A2 => n13, B1 => n573, B2 => n16, C1 
                           => n15, C2 => n607, ZN => n570);
   U519 : OAI221_X1 port map( B1 => n165, B2 => n589, C1 => n245, C2 => n608, A
                           => n609, ZN => n573);
   U520 : AOI222_X1 port map( A1 => DATA1(13), A2 => n17, B1 => DATA1(12), B2 
                           => n247, C1 => DATA1(16), C2 => n18, ZN => n609);
   U521 : AOI22_X1 port map( A1 => DATA1(16), A2 => n610, B1 => DATA2(16), B2 
                           => n611, ZN => n595);
   U522 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(16), Z => n611);
   U523 : OAI21_X1 port map( B1 => DATA2(16), B2 => n84, A => n83, ZN => n610);
   U524 : OAI211_X1 port map( C1 => n612, C2 => n123, A => n613, B => n614, ZN 
                           => OUTALU(15));
   U525 : AOI221_X1 port map( B1 => adder_out_15_port, B2 => n31, C1 => 
                           dataout_mul_15_port, C2 => n8, A => n615, ZN => n614
                           );
   U526 : NOR3_X1 port map( A1 => n113, A2 => n616, A3 => n617, ZN => n615);
   U527 : AOI22_X1 port map( A1 => DATA1(15), A2 => n618, B1 => DATA2(15), B2 
                           => n619, ZN => n613);
   U528 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(15), Z => n619);
   U529 : OAI21_X1 port map( B1 => DATA2(15), B2 => n84, A => n83, ZN => n618);
   U530 : INV_X1 port map( A => n620, ZN => n612);
   U531 : OAI22_X1 port map( A1 => n10, A2 => n581, B1 => n216, B2 => n600, ZN 
                           => n620);
   U532 : AOI221_X1 port map( B1 => n601, B2 => n221, C1 => n621, C2 => n223, A
                           => n622, ZN => n581);
   U533 : OAI222_X1 port map( A1 => n231, A2 => n603, B1 => n623, B2 => n228, 
                           C1 => n12, C2 => n547, ZN => n622);
   U534 : INV_X1 port map( A => n582, ZN => n547);
   U535 : OAI221_X1 port map( B1 => n604, B2 => n92, C1 => n624, C2 => n94, A 
                           => n625, ZN => n582);
   U536 : AOI222_X1 port map( A1 => n7, A2 => n606, B1 => n626, B2 => n375, C1 
                           => n376, C2 => n550, ZN => n625);
   U537 : INV_X1 port map( A => n585, ZN => n550);
   U538 : AOI222_X1 port map( A1 => n607, A2 => n13, B1 => n588, B2 => n16, C1 
                           => n15, C2 => n627, ZN => n585);
   U539 : OAI221_X1 port map( B1 => n165, B2 => n608, C1 => n245, C2 => n628, A
                           => n629, ZN => n588);
   U540 : AOI222_X1 port map( A1 => DATA1(12), A2 => n17, B1 => DATA1(11), B2 
                           => n247, C1 => DATA1(15), C2 => n18, ZN => n629);
   U541 : NAND2_X1 port map( A1 => n630, A2 => n631, ZN => OUTALU(14));
   U542 : AOI221_X1 port map( B1 => dataout_mul_14_port, B2 => n8, C1 => n60, 
                           C2 => n632, A => n633, ZN => n631);
   U543 : NOR3_X1 port map( A1 => n123, A2 => n600, A3 => n10, ZN => n633);
   U544 : AOI221_X1 port map( B1 => n621, B2 => n221, C1 => n634, C2 => n223, A
                           => n635, ZN => n600);
   U545 : OAI222_X1 port map( A1 => n231, A2 => n623, B1 => n636, B2 => n228, 
                           C1 => n12, C2 => n569, ZN => n635);
   U546 : INV_X1 port map( A => n601, ZN => n569);
   U547 : OAI221_X1 port map( B1 => n624, B2 => n92, C1 => n637, C2 => n94, A 
                           => n638, ZN => n601);
   U548 : AOI222_X1 port map( A1 => n7, A2 => n626, B1 => n639, B2 => n375, C1 
                           => n376, C2 => n572, ZN => n638);
   U549 : INV_X1 port map( A => n604, ZN => n572);
   U550 : AOI222_X1 port map( A1 => n627, A2 => n13, B1 => n607, B2 => n16, C1 
                           => n15, C2 => n640, ZN => n604);
   U551 : OAI221_X1 port map( B1 => n165, B2 => n628, C1 => n245, C2 => n641, A
                           => n642, ZN => n607);
   U552 : AOI222_X1 port map( A1 => DATA1(11), A2 => n17, B1 => DATA1(10), B2 
                           => n247, C1 => DATA1(14), C2 => n18, ZN => n642);
   U553 : OAI22_X1 port map( A1 => n616, A2 => n205, B1 => n643, B2 => n617, ZN
                           => n632);
   U554 : AOI21_X1 port map( B1 => adder_out_14_port, B2 => n31, A => n644, ZN 
                           => n630);
   U555 : MUX2_X1 port map( A => n645, B => n646, S => DATA2(14), Z => n644);
   U556 : NAND2_X1 port map( A1 => n647, A2 => n83, ZN => n646);
   U557 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(14), Z => n647);
   U558 : NOR2_X1 port map( A1 => n84, A2 => n608, ZN => n645);
   U559 : OAI211_X1 port map( C1 => n648, C2 => n123, A => n649, B => n650, ZN 
                           => OUTALU(13));
   U560 : AOI222_X1 port map( A1 => adder_out_13_port, A2 => n31, B1 => n60, B2
                           => n651, C1 => dataout_mul_13_port, C2 => n8, ZN => 
                           n650);
   U561 : OAI222_X1 port map( A1 => n643, A2 => n205, B1 => n652, B2 => n617, 
                           C1 => n616, C2 => n207, ZN => n651);
   U562 : INV_X1 port map( A => n653, ZN => n643);
   U563 : AOI22_X1 port map( A1 => DATA1(13), A2 => n654, B1 => DATA2(13), B2 
                           => n655, ZN => n649);
   U564 : MUX2_X1 port map( A => n337, B => n336, S => n628, Z => n655);
   U565 : OAI21_X1 port map( B1 => DATA2(13), B2 => n84, A => n83, ZN => n654);
   U566 : AOI221_X1 port map( B1 => n221, B2 => n634, C1 => n223, C2 => n656, A
                           => n657, ZN => n648);
   U567 : OAI22_X1 port map( A1 => n636, A2 => n231, B1 => n584, B2 => n12, ZN 
                           => n657);
   U568 : INV_X1 port map( A => n621, ZN => n584);
   U569 : OAI221_X1 port map( B1 => n637, B2 => n92, C1 => n658, C2 => n94, A 
                           => n659, ZN => n621);
   U570 : AOI222_X1 port map( A1 => n7, A2 => n639, B1 => n660, B2 => n375, C1 
                           => n376, C2 => n587, ZN => n659);
   U571 : INV_X1 port map( A => n624, ZN => n587);
   U572 : AOI222_X1 port map( A1 => n640, A2 => n13, B1 => n627, B2 => n16, C1 
                           => n15, C2 => n661, ZN => n624);
   U573 : OAI221_X1 port map( B1 => n165, B2 => n641, C1 => n245, C2 => n662, A
                           => n663, ZN => n627);
   U574 : AOI222_X1 port map( A1 => DATA1(10), A2 => n17, B1 => DATA1(9), B2 =>
                           n247, C1 => DATA1(13), C2 => n18, ZN => n663);
   U575 : INV_X1 port map( A => n664, ZN => n639);
   U576 : NAND2_X1 port map( A1 => n665, A2 => n666, ZN => OUTALU(12));
   U577 : AOI222_X1 port map( A1 => dataout_mul_12_port, A2 => n8, B1 => n62, 
                           B2 => n667, C1 => n60, C2 => n668, ZN => n666);
   U578 : OAI221_X1 port map( B1 => n669, B2 => n617, C1 => n616, C2 => n670, A
                           => n671, ZN => n668);
   U579 : AOI22_X1 port map( A1 => n565, A2 => n672, B1 => n564, B2 => n653, ZN
                           => n671);
   U580 : INV_X1 port map( A => n205, ZN => n565);
   U581 : INV_X1 port map( A => n673, ZN => n616);
   U582 : INV_X1 port map( A => n113, ZN => n60);
   U583 : OAI222_X1 port map( A1 => n623, A2 => n316, B1 => n603, B2 => n12, C1
                           => n636, C2 => n317, ZN => n667);
   U584 : INV_X1 port map( A => n634, ZN => n603);
   U585 : OAI221_X1 port map( B1 => n658, B2 => n92, C1 => n664, C2 => n94, A 
                           => n674, ZN => n634);
   U586 : AOI222_X1 port map( A1 => n7, A2 => n660, B1 => n69, B2 => n375, C1 
                           => n376, C2 => n606, ZN => n674);
   U587 : INV_X1 port map( A => n637, ZN => n606);
   U588 : AOI222_X1 port map( A1 => n661, A2 => n13, B1 => n640, B2 => n16, C1 
                           => n15, C2 => n675, ZN => n637);
   U589 : OAI221_X1 port map( B1 => n165, B2 => n662, C1 => n245, C2 => n676, A
                           => n677, ZN => n640);
   U590 : AOI222_X1 port map( A1 => n17, A2 => DATA1(9), B1 => DATA1(8), B2 => 
                           n247, C1 => DATA1(12), C2 => n18, ZN => n677);
   U591 : AOI21_X1 port map( B1 => adder_out_12_port, B2 => n31, A => n678, ZN 
                           => n665);
   U592 : MUX2_X1 port map( A => n679, B => n680, S => DATA2(12), Z => n678);
   U593 : NAND2_X1 port map( A1 => n681, A2 => n83, ZN => n680);
   U594 : MUX2_X1 port map( A => n85, B => n84, S => n641, Z => n681);
   U595 : NOR2_X1 port map( A1 => n84, A2 => n641, ZN => n679);
   U596 : NAND2_X1 port map( A1 => n682, A2 => n683, ZN => OUTALU(11));
   U597 : AOI221_X1 port map( B1 => dataout_mul_11_port, B2 => n8, C1 => n62, 
                           C2 => n684, A => n685, ZN => n683);
   U598 : NOR3_X1 port map( A1 => n113, A2 => n97, A3 => n96, ZN => n685);
   U599 : INV_X1 port map( A => n77, ZN => n97);
   U600 : OAI22_X1 port map( A1 => n636, A2 => n316, B1 => n623, B2 => n12, ZN 
                           => n684);
   U601 : INV_X1 port map( A => n656, ZN => n623);
   U602 : OAI221_X1 port map( B1 => n664, B2 => n92, C1 => n64, C2 => n94, A =>
                           n686, ZN => n656);
   U603 : AOI222_X1 port map( A1 => n7, A2 => n69, B1 => n71, B2 => n375, C1 =>
                           n376, C2 => n626, ZN => n686);
   U604 : INV_X1 port map( A => n658, ZN => n626);
   U605 : AOI222_X1 port map( A1 => n15, A2 => n687, B1 => n661, B2 => n16, C1 
                           => n675, C2 => n13, ZN => n658);
   U606 : OAI221_X1 port map( B1 => n165, B2 => n676, C1 => n86, C2 => n245, A 
                           => n688, ZN => n661);
   U607 : AOI222_X1 port map( A1 => DATA1(8), A2 => n17, B1 => DATA1(7), B2 => 
                           n247, C1 => DATA1(11), C2 => n18, ZN => n688);
   U608 : INV_X1 port map( A => n91, ZN => n71);
   U609 : AOI21_X1 port map( B1 => adder_out_11_port, B2 => n31, A => n689, ZN 
                           => n682);
   U610 : MUX2_X1 port map( A => n690, B => n691, S => DATA2(11), Z => n689);
   U611 : NAND2_X1 port map( A1 => n692, A2 => n83, ZN => n691);
   U612 : MUX2_X1 port map( A => n84, B => n85, S => DATA1(11), Z => n692);
   U613 : NOR2_X1 port map( A1 => n84, A2 => n662, ZN => n690);
   U614 : OAI211_X1 port map( C1 => n693, C2 => n113, A => n694, B => n695, ZN 
                           => OUTALU(10));
   U615 : AOI221_X1 port map( B1 => adder_out_10_port, B2 => n31, C1 => 
                           dataout_mul_10_port, C2 => n8, A => n696, ZN => n695
                           );
   U616 : NOR3_X1 port map( A1 => n123, A2 => n636, A3 => n12, ZN => n696);
   U617 : AOI221_X1 port map( B1 => n660, B2 => n68, C1 => n69, C2 => n70, A =>
                           n697, ZN => n636);
   U618 : OAI222_X1 port map( A1 => n2, A2 => n91, B1 => n66, B2 => n237, C1 =>
                           n65, C2 => n664, ZN => n697);
   U619 : AOI222_X1 port map( A1 => n15, A2 => n698, B1 => n687, B2 => n13, C1 
                           => n675, C2 => n16, ZN => n664);
   U620 : OAI221_X1 port map( B1 => n86, B2 => n165, C1 => n245, C2 => n106, A 
                           => n699, ZN => n675);
   U621 : AOI222_X1 port map( A1 => DATA1(7), A2 => n17, B1 => DATA1(6), B2 => 
                           n247, C1 => DATA1(10), C2 => n18, ZN => n699);
   U622 : AOI222_X1 port map( A1 => n15, A2 => n138, B1 => n140, B2 => n13, C1 
                           => n700, C2 => n16, ZN => n66);
   U623 : OAI221_X1 port map( B1 => n165, B2 => n164, C1 => n245, C2 => n166, A
                           => n701, ZN => n138);
   U624 : AOI222_X1 port map( A1 => DATA1(1), A2 => n17, B1 => DATA1(0), B2 => 
                           n247, C1 => DATA1(4), C2 => n18, ZN => n701);
   U625 : AOI222_X1 port map( A1 => n702, A2 => n16, B1 => n15, B2 => n140, C1 
                           => n700, C2 => n13, ZN => n91);
   U626 : OAI221_X1 port map( B1 => n165, B2 => n156, C1 => n245, C2 => n164, A
                           => n703, ZN => n140);
   U627 : AOI222_X1 port map( A1 => DATA1(2), A2 => n17, B1 => DATA1(1), B2 => 
                           n247, C1 => DATA1(5), C2 => n18, ZN => n703);
   U628 : INV_X1 port map( A => n93, ZN => n69);
   U629 : AOI222_X1 port map( A1 => n15, A2 => n700, B1 => n702, B2 => n13, C1 
                           => n698, C2 => n16, ZN => n93);
   U630 : OAI221_X1 port map( B1 => n165, B2 => n145, C1 => n245, C2 => n156, A
                           => n704, ZN => n700);
   U631 : AOI222_X1 port map( A1 => DATA1(3), A2 => n17, B1 => DATA1(2), B2 => 
                           n247, C1 => DATA1(6), C2 => n18, ZN => n704);
   U632 : INV_X1 port map( A => n64, ZN => n660);
   U633 : AOI222_X1 port map( A1 => n687, A2 => n16, B1 => n15, B2 => n702, C1 
                           => n698, C2 => n13, ZN => n64);
   U634 : OAI221_X1 port map( B1 => n165, B2 => n118, C1 => n245, C2 => n130, A
                           => n705, ZN => n698);
   U635 : AOI222_X1 port map( A1 => DATA1(5), A2 => n17, B1 => DATA1(4), B2 => 
                           n247, C1 => DATA1(8), C2 => n18, ZN => n705);
   U636 : OAI221_X1 port map( B1 => n165, B2 => n130, C1 => n245, C2 => n145, A
                           => n706, ZN => n702);
   U637 : AOI222_X1 port map( A1 => DATA1(4), A2 => n17, B1 => DATA1(3), B2 => 
                           n247, C1 => DATA1(7), C2 => n18, ZN => n706);
   U638 : OAI221_X1 port map( B1 => n165, B2 => n106, C1 => n245, C2 => n118, A
                           => n707, ZN => n687);
   U639 : AOI222_X1 port map( A1 => DATA1(6), A2 => n17, B1 => DATA1(5), B2 => 
                           n247, C1 => DATA1(9), C2 => n18, ZN => n707);
   U640 : INV_X1 port map( A => n62, ZN => n123);
   U641 : AOI22_X1 port map( A1 => DATA1(10), A2 => n708, B1 => DATA2(10), B2 
                           => n709, ZN => n694);
   U642 : MUX2_X1 port map( A => n337, B => n336, S => n676, Z => n709);
   U643 : OAI21_X1 port map( B1 => DATA2(10), B2 => n84, A => n83, ZN => n708);
   U644 : AOI22_X1 port map( A1 => n76, A2 => n73, B1 => n74, B2 => n77, ZN => 
                           n693);
   U645 : NAND4_X1 port map( A1 => n710, A2 => n711, A3 => n712, A4 => n713, ZN
                           => OUTALU(0));
   U646 : AOI221_X1 port map( B1 => n714, B2 => n62, C1 => DATA2(0), C2 => n715
                           , A => n716, ZN => n713);
   U647 : OAI21_X1 port map( B1 => n717, B2 => n294, A => n718, ZN => n716);
   U648 : NAND3_X1 port map( A1 => FUNC(0), A2 => n719, A3 => n720, ZN => n718)
                           ;
   U649 : MUX2_X1 port map( A => n721, B => n722, S => FUNC(2), Z => n720);
   U650 : AND2_X1 port map( A1 => N2515, A2 => n723, ZN => n722);
   U651 : MUX2_X1 port map( A => N2513, B => N2514, S => FUNC(3), Z => n721);
   U652 : AOI21_X1 port map( B1 => n336, B2 => n724, A => n725, ZN => n717);
   U653 : INV_X1 port map( A => n83, ZN => n725);
   U654 : MUX2_X1 port map( A => n336, B => n337, S => DATA1(0), Z => n715);
   U655 : INV_X1 port map( A => n85, ZN => n337);
   U656 : NAND3_X1 port map( A1 => FUNC(2), A2 => n728, A3 => FUNC(3), ZN => 
                           n85);
   U657 : INV_X1 port map( A => n84, ZN => n336);
   U658 : NAND3_X1 port map( A1 => FUNC(2), A2 => n723, A3 => n727, ZN => n252)
                           ;
   U659 : AOI22_X1 port map( A1 => dataout_mul_0_port, A2 => n8, B1 => 
                           adder_out_0_port, B2 => n31, ZN => n712);
   U660 : INV_X1 port map( A => n20, ZN => n730);
   U661 : NAND4_X1 port map( A1 => n18, A2 => n731, A3 => n732, A4 => n733, ZN 
                           => n20);
   U662 : NOR4_X1 port map( A1 => n734, A2 => DATA2(14), A3 => DATA2(6), A4 => 
                           DATA2(15), ZN => n733);
   U663 : OR3_X1 port map( A1 => DATA2(8), A2 => DATA2(9), A3 => DATA2(7), ZN 
                           => n734);
   U664 : NOR3_X1 port map( A1 => DATA2(11), A2 => DATA2(13), A3 => DATA2(12), 
                           ZN => n732);
   U665 : INV_X1 port map( A => DATA2(10), ZN => n731);
   U666 : INV_X1 port map( A => n19, ZN => n1034);
   U667 : NAND4_X1 port map( A1 => n735, A2 => n736, A3 => n737, A4 => n738, ZN
                           => n19);
   U668 : NOR4_X1 port map( A1 => DATA1(9), A2 => DATA1(8), A3 => DATA1(7), A4 
                           => DATA1(6), ZN => n738);
   U669 : NOR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(3), A4 
                           => DATA1(2), ZN => n737);
   U670 : NOR4_X1 port map( A1 => DATA1(1), A2 => DATA1(15), A3 => DATA1(14), 
                           A4 => DATA1(13), ZN => n736);
   U671 : NOR4_X1 port map( A1 => DATA1(12), A2 => DATA1(11), A3 => DATA1(10), 
                           A4 => DATA1(0), ZN => n735);
   U672 : NAND4_X1 port map( A1 => n739, A2 => n531, A3 => n729, A4 => n740, ZN
                           => n711);
   U673 : OAI221_X1 port map( B1 => n289, B2 => n150, C1 => n161, C2 => n162, A
                           => n741, ZN => n531);
   U674 : AOI222_X1 port map( A1 => n190, A2 => n163, B1 => n186, B2 => n293, 
                           C1 => n188, C2 => n742, ZN => n741);
   U675 : OAI222_X1 port map( A1 => n743, A2 => n111, B1 => n192, B2 => n112, 
                           C1 => n124, C2 => n125, ZN => n293);
   U676 : AOI221_X1 port map( B1 => n101, B2 => n74, C1 => n75, C2 => n78, A =>
                           n744, ZN => n112);
   U677 : INV_X1 port map( A => n745, ZN => n744);
   U678 : AOI222_X1 port map( A1 => n199, A2 => n73, B1 => n201, B2 => n77, C1 
                           => n76, C2 => n746, ZN => n745);
   U679 : OAI221_X1 port map( B1 => n669, B2 => n205, C1 => n652, C2 => n207, A
                           => n747, ZN => n77);
   U680 : AOI222_X1 port map( A1 => n209, A2 => n653, B1 => n214, B2 => n673, 
                           C1 => n212, C2 => n748, ZN => n747);
   U681 : OAI222_X1 port map( A1 => n219, A2 => n579, B1 => n749, B2 => n10, C1
                           => n599, C2 => n216, ZN => n673);
   U682 : AOI221_X1 port map( B1 => n750, B2 => n221, C1 => n751, C2 => n223, A
                           => n752, ZN => n579);
   U683 : OAI222_X1 port map( A1 => n231, A2 => n514, B1 => n494, B2 => n228, 
                           C1 => n12, C2 => n753, ZN => n752);
   U684 : AOI221_X1 port map( B1 => n474, B2 => n68, C1 => n754, C2 => n70, A 
                           => n755, ZN => n494);
   U685 : OAI222_X1 port map( A1 => n2, A2 => n431, B1 => n409, B2 => n237, C1 
                           => n65, C2 => n756, ZN => n755);
   U686 : AOI222_X1 port map( A1 => n757, A2 => n16, B1 => n15, B2 => n359, C1 
                           => n384, C2 => n13, ZN => n409);
   U687 : OAI221_X1 port map( B1 => n55, B2 => n165, C1 => n56, C2 => n245, A 
                           => n758, ZN => n359);
   U688 : AOI222_X1 port map( A1 => DATA1(30), A2 => n17, B1 => DATA1(31), B2 
                           => n247, C1 => DATA1(27), C2 => n18, ZN => n758);
   U689 : INV_X1 port map( A => DATA1(29), ZN => n56);
   U690 : INV_X1 port map( A => n672, ZN => n652);
   U691 : INV_X1 port map( A => n181, ZN => n162);
   U692 : INV_X1 port map( A => n292, ZN => n161);
   U693 : INV_X1 port map( A => n759, ZN => n289);
   U694 : INV_X1 port map( A => n760, ZN => n710);
   U695 : AOI21_X1 port map( B1 => n761, B2 => n762, A => n113, ZN => n760);
   U696 : NAND2_X1 port map( A1 => n739, A2 => n250, ZN => n113);
   U697 : INV_X1 port map( A => n729, ZN => n250);
   U698 : OAI21_X1 port map( B1 => n763, B2 => n764, A => n740, ZN => n729);
   U699 : INV_X1 port map( A => DATA2(5), ZN => n740);
   U700 : AND3_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n727, ZN => 
                           n739);
   U701 : NOR2_X1 port map( A1 => n719, A2 => FUNC(0), ZN => n727);
   U702 : INV_X1 port map( A => FUNC(1), ZN => n719);
   U703 : AOI22_X1 port map( A1 => n759, A2 => n181, B1 => n742, B2 => n179, ZN
                           => n762);
   U704 : INV_X1 port map( A => n150, ZN => n179);
   U705 : NAND2_X1 port map( A1 => n135, A2 => n765, ZN => n150);
   U706 : OAI222_X1 port map( A1 => n766, A2 => n125, B1 => n767, B2 => n111, 
                           C1 => n192, C2 => n768, ZN => n742);
   U707 : NOR2_X1 port map( A1 => n765, A2 => n769, ZN => n181);
   U708 : OAI222_X1 port map( A1 => n192, A2 => n770, B1 => n768, B2 => n125, 
                           C1 => n766, C2 => n111, ZN => n759);
   U709 : AOI222_X1 port map( A1 => n163, A2 => n186, B1 => n771, B2 => n188, 
                           C1 => n292, C2 => n190, ZN => n761);
   U710 : INV_X1 port map( A => n290, ZN => n190);
   U711 : NAND2_X1 port map( A1 => n769, A2 => n772, ZN => n290);
   U712 : OAI21_X1 port map( B1 => n773, B2 => n763, A => n772, ZN => n769);
   U713 : OAI222_X1 port map( A1 => n770, A2 => n125, B1 => n192, B2 => n743, 
                           C1 => n768, C2 => n111, ZN => n292);
   U714 : AOI221_X1 port map( B1 => n774, B2 => n74, C1 => n775, C2 => n78, A 
                           => n776, ZN => n768);
   U715 : INV_X1 port map( A => n777, ZN => n776);
   U716 : AOI222_X1 port map( A1 => n199, A2 => n778, B1 => n201, B2 => n746, 
                           C1 => n76, C2 => n779, ZN => n777);
   U717 : INV_X1 port map( A => n135, ZN => n188);
   U718 : OAI21_X1 port map( B1 => n764, B2 => n780, A => n765, ZN => n135);
   U719 : OAI222_X1 port map( A1 => n766, A2 => n192, B1 => n111, B2 => n781, 
                           C1 => n125, C2 => n767, ZN => n771);
   U720 : AOI221_X1 port map( B1 => n782, B2 => n74, C1 => n779, C2 => n78, A 
                           => n783, ZN => n767);
   U721 : INV_X1 port map( A => n784, ZN => n783);
   U722 : AOI222_X1 port map( A1 => n199, A2 => n774, B1 => n201, B2 => n775, 
                           C1 => n76, C2 => n785, ZN => n784);
   U723 : AOI221_X1 port map( B1 => n785, B2 => n74, C1 => n782, C2 => n78, A 
                           => n786, ZN => n781);
   U724 : INV_X1 port map( A => n787, ZN => n786);
   U725 : AOI222_X1 port map( A1 => n199, A2 => n779, B1 => n201, B2 => n774, 
                           C1 => n76, C2 => n788, ZN => n787);
   U726 : OAI221_X1 port map( B1 => n789, B2 => n205, C1 => n790, C2 => n207, A
                           => n791, ZN => n788);
   U727 : AOI222_X1 port map( A1 => n209, A2 => n792, B1 => n793, B2 => n212, 
                           C1 => n794, C2 => n214, ZN => n791);
   U728 : OAI222_X1 port map( A1 => n795, A2 => n216, B1 => n796, B2 => n10, C1
                           => n219, C2 => n797, ZN => n793);
   U729 : INV_X1 port map( A => n798, ZN => n796);
   U730 : OAI221_X1 port map( B1 => n316, B2 => n799, C1 => n317, C2 => n800, A
                           => n801, ZN => n798);
   U731 : AOI222_X1 port map( A1 => n802, A2 => n11, B1 => n274, B2 => n803, C1
                           => n804, C2 => n271, ZN => n801);
   U732 : OAI221_X1 port map( B1 => n92, B2 => n805, C1 => n94, C2 => n806, A 
                           => n807, ZN => n802);
   U733 : INV_X1 port map( A => n808, ZN => n807);
   U734 : OAI222_X1 port map( A1 => n237, A2 => n809, B1 => n810, B2 => n65, C1
                           => n811, C2 => n2, ZN => n808);
   U735 : AOI222_X1 port map( A1 => n812, A2 => n15, B1 => n16, B2 => n813, C1 
                           => n13, C2 => n814, ZN => n810);
   U736 : OAI221_X1 port map( B1 => n165, B2 => n295, C1 => n245, C2 => n166, A
                           => n815, ZN => n813);
   U737 : AOI221_X1 port map( B1 => DATA1(3), B2 => n17, C1 => DATA1(4), C2 => 
                           n247, A => n714, ZN => n815);
   U738 : NOR2_X1 port map( A1 => n294, A2 => n3, ZN => n714);
   U739 : INV_X1 port map( A => DATA1(0), ZN => n294);
   U740 : INV_X1 port map( A => DATA1(1), ZN => n295);
   U741 : INV_X1 port map( A => n223, ZN => n317);
   U742 : INV_X1 port map( A => n816, ZN => n789);
   U743 : OAI221_X1 port map( B1 => n790, B2 => n205, C1 => n817, C2 => n207, A
                           => n818, ZN => n785);
   U744 : AOI222_X1 port map( A1 => n209, A2 => n794, B1 => n819, B2 => n214, 
                           C1 => n816, C2 => n212, ZN => n818);
   U745 : OAI222_X1 port map( A1 => n219, A2 => n820, B1 => n795, B2 => n10, C1
                           => n797, C2 => n216, ZN => n816);
   U746 : AOI221_X1 port map( B1 => n821, B2 => n221, C1 => n804, C2 => n223, A
                           => n822, ZN => n795);
   U747 : OAI222_X1 port map( A1 => n231, A2 => n823, B1 => n824, B2 => n228, 
                           C1 => n12, C2 => n799, ZN => n822);
   U748 : AOI221_X1 port map( B1 => n825, B2 => n68, C1 => n826, C2 => n70, A 
                           => n827, ZN => n799);
   U749 : OAI222_X1 port map( A1 => n2, A2 => n809, B1 => n828, B2 => n237, C1 
                           => n65, C2 => n805, ZN => n827);
   U750 : AOI222_X1 port map( A1 => n15, A2 => n829, B1 => n814, B2 => n16, C1 
                           => n812, C2 => n13, ZN => n805);
   U751 : OAI221_X1 port map( B1 => n165, B2 => n166, C1 => n245, C2 => n164, A
                           => n830, ZN => n814);
   U752 : AOI222_X1 port map( A1 => DATA1(4), A2 => n17, B1 => DATA1(5), B2 => 
                           n247, C1 => DATA1(1), C2 => n18, ZN => n830);
   U753 : INV_X1 port map( A => DATA1(2), ZN => n166);
   U754 : INV_X1 port map( A => n806, ZN => n825);
   U755 : INV_X1 port map( A => n800, ZN => n821);
   U756 : INV_X1 port map( A => n831, ZN => n790);
   U757 : AOI221_X1 port map( B1 => n779, B2 => n74, C1 => n774, C2 => n78, A 
                           => n832, ZN => n766);
   U758 : INV_X1 port map( A => n833, ZN => n832);
   U759 : AOI222_X1 port map( A1 => n199, A2 => n775, B1 => n201, B2 => n778, 
                           C1 => n76, C2 => n782, ZN => n833);
   U760 : OAI221_X1 port map( B1 => n817, B2 => n205, C1 => n834, C2 => n207, A
                           => n835, ZN => n782);
   U761 : AOI222_X1 port map( A1 => n209, A2 => n819, B1 => n836, B2 => n214, 
                           C1 => n831, C2 => n212, ZN => n835);
   U762 : OAI222_X1 port map( A1 => n219, A2 => n837, B1 => n820, B2 => n216, 
                           C1 => n797, C2 => n10, ZN => n831);
   U763 : AOI221_X1 port map( B1 => n804, B2 => n221, C1 => n803, C2 => n223, A
                           => n838, ZN => n797);
   U764 : OAI222_X1 port map( A1 => n231, A2 => n824, B1 => n839, B2 => n228, 
                           C1 => n12, C2 => n800, ZN => n838);
   U765 : AOI221_X1 port map( B1 => n826, B2 => n68, C1 => n840, C2 => n70, A 
                           => n841, ZN => n800);
   U766 : OAI222_X1 port map( A1 => n2, A2 => n828, B1 => n237, B2 => n842, C1 
                           => n65, C2 => n806, ZN => n841);
   U767 : AOI222_X1 port map( A1 => n15, A2 => n843, B1 => n829, B2 => n13, C1 
                           => n812, C2 => n16, ZN => n806);
   U768 : OAI221_X1 port map( B1 => n165, B2 => n164, C1 => n245, C2 => n156, A
                           => n844, ZN => n812);
   U769 : AOI222_X1 port map( A1 => DATA1(5), A2 => n17, B1 => DATA1(6), B2 => 
                           n247, C1 => DATA1(2), C2 => n18, ZN => n844);
   U770 : INV_X1 port map( A => DATA1(3), ZN => n164);
   U771 : INV_X1 port map( A => n792, ZN => n817);
   U772 : OAI221_X1 port map( B1 => n834, B2 => n205, C1 => n845, C2 => n207, A
                           => n846, ZN => n779);
   U773 : AOI222_X1 port map( A1 => n209, A2 => n836, B1 => n847, B2 => n214, 
                           C1 => n792, C2 => n212, ZN => n846);
   U774 : OAI222_X1 port map( A1 => n820, A2 => n10, B1 => n219, B2 => n848, C1
                           => n837, C2 => n216, ZN => n792);
   U775 : AOI221_X1 port map( B1 => n803, B2 => n221, C1 => n849, C2 => n223, A
                           => n850, ZN => n820);
   U776 : INV_X1 port map( A => n851, ZN => n850);
   U777 : AOI222_X1 port map( A1 => n271, A2 => n852, B1 => n853, B2 => n274, 
                           C1 => n11, C2 => n804, ZN => n851);
   U778 : OAI221_X1 port map( B1 => n809, B2 => n92, C1 => n828, C2 => n94, A 
                           => n854, ZN => n804);
   U779 : AOI222_X1 port map( A1 => n7, A2 => n855, B1 => n375, B2 => n856, C1 
                           => n376, C2 => n826, ZN => n854);
   U780 : INV_X1 port map( A => n811, ZN => n826);
   U781 : AOI222_X1 port map( A1 => n829, A2 => n16, B1 => n15, B2 => n857, C1 
                           => n843, C2 => n13, ZN => n811);
   U782 : OAI221_X1 port map( B1 => n165, B2 => n156, C1 => n245, C2 => n145, A
                           => n858, ZN => n829);
   U783 : AOI222_X1 port map( A1 => DATA1(6), A2 => n17, B1 => DATA1(7), B2 => 
                           n247, C1 => DATA1(3), C2 => n18, ZN => n858);
   U784 : INV_X1 port map( A => DATA1(4), ZN => n156);
   U785 : INV_X1 port map( A => n231, ZN => n271);
   U786 : INV_X1 port map( A => n794, ZN => n834);
   U787 : INV_X1 port map( A => n772, ZN => n186);
   U788 : NAND2_X1 port map( A1 => n859, A2 => n860, ZN => n772);
   U789 : OAI222_X1 port map( A1 => n192, A2 => n124, B1 => n743, B2 => n125, 
                           C1 => n770, C2 => n111, ZN => n163);
   U790 : AOI221_X1 port map( B1 => n775, B2 => n74, C1 => n778, C2 => n78, A 
                           => n861, ZN => n770);
   U791 : INV_X1 port map( A => n862, ZN => n861);
   U792 : AOI222_X1 port map( A1 => n199, A2 => n746, B1 => n201, B2 => n101, 
                           C1 => n76, C2 => n774, ZN => n862);
   U793 : OAI221_X1 port map( B1 => n845, B2 => n205, C1 => n863, C2 => n207, A
                           => n864, ZN => n774);
   U794 : AOI222_X1 port map( A1 => n209, A2 => n847, B1 => n865, B2 => n214, 
                           C1 => n794, C2 => n212, ZN => n864);
   U795 : OAI222_X1 port map( A1 => n219, A2 => n866, B1 => n848, B2 => n216, 
                           C1 => n837, C2 => n10, ZN => n794);
   U796 : AOI221_X1 port map( B1 => n849, B2 => n221, C1 => n852, C2 => n223, A
                           => n867, ZN => n837);
   U797 : OAI222_X1 port map( A1 => n231, A2 => n868, B1 => n869, B2 => n228, 
                           C1 => n12, C2 => n823, ZN => n867);
   U798 : INV_X1 port map( A => n803, ZN => n823);
   U799 : OAI221_X1 port map( B1 => n828, B2 => n92, C1 => n842, C2 => n94, A 
                           => n870, ZN => n803);
   U800 : AOI222_X1 port map( A1 => n7, A2 => n856, B1 => n375, B2 => n871, C1 
                           => n376, C2 => n840, ZN => n870);
   U801 : INV_X1 port map( A => n809, ZN => n840);
   U802 : AOI222_X1 port map( A1 => n15, A2 => n872, B1 => n857, B2 => n13, C1 
                           => n843, C2 => n16, ZN => n809);
   U803 : OAI221_X1 port map( B1 => n165, B2 => n145, C1 => n245, C2 => n130, A
                           => n873, ZN => n843);
   U804 : AOI222_X1 port map( A1 => DATA1(7), A2 => n17, B1 => DATA1(8), B2 => 
                           n247, C1 => DATA1(4), C2 => n18, ZN => n873);
   U805 : INV_X1 port map( A => DATA1(5), ZN => n145);
   U806 : INV_X1 port map( A => n824, ZN => n849);
   U807 : INV_X1 port map( A => n819, ZN => n845);
   U808 : NAND2_X1 port map( A1 => n192, A2 => n111, ZN => n125);
   U809 : AOI221_X1 port map( B1 => n778, B2 => n74, C1 => n746, C2 => n78, A 
                           => n874, ZN => n743);
   U810 : INV_X1 port map( A => n875, ZN => n874);
   U811 : AOI222_X1 port map( A1 => n199, A2 => n101, B1 => n201, B2 => n75, C1
                           => n76, C2 => n775, ZN => n875);
   U812 : OAI221_X1 port map( B1 => n863, B2 => n205, C1 => n876, C2 => n207, A
                           => n877, ZN => n775);
   U813 : AOI222_X1 port map( A1 => n209, A2 => n865, B1 => n878, B2 => n214, 
                           C1 => n819, C2 => n212, ZN => n877);
   U814 : OAI222_X1 port map( A1 => n848, A2 => n10, B1 => n219, B2 => n879, C1
                           => n866, C2 => n216, ZN => n819);
   U815 : AOI221_X1 port map( B1 => n852, B2 => n221, C1 => n853, C2 => n223, A
                           => n880, ZN => n848);
   U816 : OAI222_X1 port map( A1 => n231, A2 => n869, B1 => n881, B2 => n228, 
                           C1 => n12, C2 => n824, ZN => n880);
   U817 : AOI221_X1 port map( B1 => n855, B2 => n68, C1 => n856, C2 => n70, A 
                           => n882, ZN => n824);
   U818 : OAI222_X1 port map( A1 => n2, A2 => n883, B1 => n237, B2 => n884, C1 
                           => n65, C2 => n828, ZN => n882);
   U819 : AOI222_X1 port map( A1 => n857, A2 => n16, B1 => n15, B2 => n885, C1 
                           => n872, C2 => n13, ZN => n828);
   U820 : OAI221_X1 port map( B1 => n165, B2 => n130, C1 => n245, C2 => n118, A
                           => n886, ZN => n857);
   U821 : AOI222_X1 port map( A1 => DATA1(8), A2 => n17, B1 => DATA1(9), B2 => 
                           n247, C1 => DATA1(5), C2 => n18, ZN => n886);
   U822 : INV_X1 port map( A => DATA1(6), ZN => n130);
   U823 : INV_X1 port map( A => n842, ZN => n855);
   U824 : INV_X1 port map( A => n839, ZN => n852);
   U825 : INV_X1 port map( A => n836, ZN => n863);
   U826 : AOI221_X1 port map( B1 => n746, B2 => n74, C1 => n101, C2 => n78, A 
                           => n887, ZN => n124);
   U827 : INV_X1 port map( A => n888, ZN => n887);
   U828 : AOI222_X1 port map( A1 => n199, A2 => n75, B1 => n201, B2 => n73, C1 
                           => n76, C2 => n778, ZN => n888);
   U829 : OAI221_X1 port map( B1 => n876, B2 => n205, C1 => n889, C2 => n207, A
                           => n890, ZN => n778);
   U830 : AOI222_X1 port map( A1 => n209, A2 => n878, B1 => n214, B2 => n891, 
                           C1 => n836, C2 => n212, ZN => n890);
   U831 : OAI222_X1 port map( A1 => n219, A2 => n892, B1 => n879, B2 => n216, 
                           C1 => n866, C2 => n10, ZN => n836);
   U832 : AOI221_X1 port map( B1 => n853, B2 => n221, C1 => n893, C2 => n223, A
                           => n894, ZN => n866);
   U833 : OAI222_X1 port map( A1 => n231, A2 => n881, B1 => n228, B2 => n895, 
                           C1 => n12, C2 => n839, ZN => n894);
   U834 : AOI221_X1 port map( B1 => n856, B2 => n68, C1 => n871, C2 => n70, A 
                           => n896, ZN => n839);
   U835 : OAI222_X1 port map( A1 => n2, A2 => n884, B1 => n237, B2 => n897, C1 
                           => n65, C2 => n842, ZN => n896);
   U836 : AOI222_X1 port map( A1 => n15, A2 => n898, B1 => n872, B2 => n16, C1 
                           => n885, C2 => n13, ZN => n842);
   U837 : OAI221_X1 port map( B1 => n165, B2 => n118, C1 => n245, C2 => n106, A
                           => n899, ZN => n872);
   U838 : AOI222_X1 port map( A1 => n17, A2 => DATA1(9), B1 => DATA1(10), B2 =>
                           n247, C1 => DATA1(6), C2 => n18, ZN => n899);
   U839 : INV_X1 port map( A => DATA1(7), ZN => n118);
   U840 : INV_X1 port map( A => n847, ZN => n876);
   U841 : INV_X1 port map( A => n96, ZN => n76);
   U842 : OAI221_X1 port map( B1 => n900, B2 => n205, C1 => n669, C2 => n207, A
                           => n901, ZN => n73);
   U843 : AOI222_X1 port map( A1 => n209, A2 => n672, B1 => n214, B2 => n653, 
                           C1 => n212, C2 => n891, ZN => n901);
   U844 : OAI222_X1 port map( A1 => n219, A2 => n599, B1 => n902, B2 => n10, C1
                           => n749, C2 => n216, ZN => n653);
   U845 : AOI221_X1 port map( B1 => n903, B2 => n221, C1 => n750, C2 => n223, A
                           => n904, ZN => n599);
   U846 : OAI222_X1 port map( A1 => n231, A2 => n539, B1 => n514, B2 => n228, 
                           C1 => n12, C2 => n905, ZN => n904);
   U847 : AOI221_X1 port map( B1 => n906, B2 => n68, C1 => n474, C2 => n70, A 
                           => n907, ZN => n514);
   U848 : OAI222_X1 port map( A1 => n2, A2 => n453, B1 => n431, B2 => n237, C1 
                           => n65, C2 => n908, ZN => n907);
   U849 : AOI222_X1 port map( A1 => n15, A2 => n384, B1 => n757, B2 => n13, C1 
                           => n909, C2 => n16, ZN => n431);
   U850 : OAI221_X1 port map( B1 => n165, B2 => n54, C1 => n55, C2 => n245, A 
                           => n910, ZN => n384);
   U851 : AOI222_X1 port map( A1 => n17, A2 => DATA1(29), B1 => DATA1(30), B2 
                           => n247, C1 => DATA1(26), C2 => n18, ZN => n910);
   U852 : INV_X1 port map( A => DATA1(28), ZN => n55);
   U853 : INV_X1 port map( A => n911, ZN => n669);
   U854 : OAI221_X1 port map( B1 => n912, B2 => n205, C1 => n900, C2 => n207, A
                           => n913, ZN => n75);
   U855 : AOI222_X1 port map( A1 => n209, A2 => n911, B1 => n214, B2 => n672, 
                           C1 => n878, C2 => n212, ZN => n913);
   U856 : OAI222_X1 port map( A1 => n914, A2 => n10, B1 => n219, B2 => n749, C1
                           => n902, C2 => n216, ZN => n672);
   U857 : AOI221_X1 port map( B1 => n915, B2 => n221, C1 => n903, C2 => n223, A
                           => n916, ZN => n749);
   U858 : OAI222_X1 port map( A1 => n231, A2 => n559, B1 => n539, B2 => n228, 
                           C1 => n12, C2 => n917, ZN => n916);
   U859 : INV_X1 port map( A => n751, ZN => n539);
   U860 : OAI221_X1 port map( B1 => n908, B2 => n92, C1 => n756, C2 => n94, A 
                           => n918, ZN => n751);
   U861 : AOI222_X1 port map( A1 => n7, A2 => n474, B1 => n754, B2 => n375, C1 
                           => n376, C2 => n919, ZN => n918);
   U862 : INV_X1 port map( A => n453, ZN => n754);
   U863 : AOI222_X1 port map( A1 => n920, A2 => n16, B1 => n15, B2 => n757, C1 
                           => n909, C2 => n13, ZN => n453);
   U864 : OAI221_X1 port map( B1 => n165, B2 => n53, C1 => n245, C2 => n54, A 
                           => n921, ZN => n757);
   U865 : AOI222_X1 port map( A1 => DATA1(28), A2 => n17, B1 => DATA1(29), B2 
                           => n247, C1 => DATA1(25), C2 => n18, ZN => n921);
   U866 : INV_X1 port map( A => DATA1(27), ZN => n54);
   U867 : INV_X1 port map( A => n748, ZN => n900);
   U868 : INV_X1 port map( A => n99, ZN => n199);
   U869 : NAND2_X1 port map( A1 => n922, A2 => n923, ZN => n99);
   U870 : OAI21_X1 port map( B1 => n925, B2 => n763, A => n923, ZN => n922);
   U871 : OAI221_X1 port map( B1 => n926, B2 => n205, C1 => n912, C2 => n207, A
                           => n927, ZN => n101);
   U872 : AOI222_X1 port map( A1 => n209, A2 => n748, B1 => n214, B2 => n911, 
                           C1 => n865, C2 => n212, ZN => n927);
   U873 : OAI222_X1 port map( A1 => n219, A2 => n902, B1 => n914, B2 => n216, 
                           C1 => n928, C2 => n10, ZN => n911);
   U874 : AOI221_X1 port map( B1 => n929, B2 => n221, C1 => n915, C2 => n223, A
                           => n930, ZN => n902);
   U875 : OAI222_X1 port map( A1 => n231, A2 => n753, B1 => n559, B2 => n228, 
                           C1 => n12, C2 => n931, ZN => n930);
   U876 : INV_X1 port map( A => n750, ZN => n559);
   U877 : OAI221_X1 port map( B1 => n932, B2 => n92, C1 => n908, C2 => n94, A 
                           => n933, ZN => n750);
   U878 : AOI222_X1 port map( A1 => n7, A2 => n906, B1 => n474, B2 => n375, C1 
                           => n376, C2 => n934, ZN => n933);
   U879 : INV_X1 port map( A => n935, ZN => n474);
   U880 : AOI222_X1 port map( A1 => n15, A2 => n909, B1 => n920, B2 => n13, C1 
                           => n936, C2 => n16, ZN => n935);
   U881 : OAI221_X1 port map( B1 => n52, B2 => n165, C1 => n53, C2 => n245, A 
                           => n937, ZN => n909);
   U882 : AOI222_X1 port map( A1 => DATA1(27), A2 => n17, B1 => DATA1(28), B2 
                           => n247, C1 => DATA1(24), C2 => n18, ZN => n937);
   U883 : INV_X1 port map( A => DATA1(26), ZN => n53);
   U884 : INV_X1 port map( A => n891, ZN => n912);
   U885 : AND2_X1 port map( A1 => n924, A2 => n96, ZN => n74);
   U886 : NAND2_X1 port map( A1 => n924, A2 => n763, ZN => n96);
   U887 : NAND2_X1 port map( A1 => DATA2(0), A2 => n860, ZN => n763);
   U888 : AOI21_X1 port map( B1 => DATA2(1), B2 => n860, A => n201, ZN => n924)
                           ;
   U889 : OAI221_X1 port map( B1 => n889, B2 => n205, C1 => n926, C2 => n207, A
                           => n938, ZN => n746);
   U890 : AOI222_X1 port map( A1 => n209, A2 => n891, B1 => n214, B2 => n748, 
                           C1 => n847, C2 => n212, ZN => n938);
   U891 : OAI222_X1 port map( A1 => n879, A2 => n10, B1 => n219, B2 => n939, C1
                           => n892, C2 => n216, ZN => n847);
   U892 : AOI221_X1 port map( B1 => n893, B2 => n221, C1 => n940, C2 => n223, A
                           => n941, ZN => n879);
   U893 : OAI222_X1 port map( A1 => n231, A2 => n895, B1 => n228, B2 => n942, 
                           C1 => n12, C2 => n868, ZN => n941);
   U894 : INV_X1 port map( A => n853, ZN => n868);
   U895 : OAI221_X1 port map( B1 => n883, B2 => n92, C1 => n884, C2 => n94, A 
                           => n943, ZN => n853);
   U896 : AOI222_X1 port map( A1 => n7, A2 => n944, B1 => n375, B2 => n945, C1 
                           => n376, C2 => n856, ZN => n943);
   U897 : INV_X1 port map( A => n946, ZN => n856);
   U898 : AOI222_X1 port map( A1 => n15, A2 => n947, B1 => n885, B2 => n16, C1 
                           => n898, C2 => n13, ZN => n946);
   U899 : OAI221_X1 port map( B1 => n165, B2 => n106, C1 => n86, C2 => n245, A 
                           => n948, ZN => n885);
   U900 : AOI222_X1 port map( A1 => DATA1(10), A2 => n17, B1 => DATA1(11), B2 
                           => n247, C1 => DATA1(7), C2 => n18, ZN => n948);
   U901 : INV_X1 port map( A => DATA1(8), ZN => n106);
   U902 : OAI222_X1 port map( A1 => n949, A2 => n10, B1 => n219, B2 => n914, C1
                           => n928, C2 => n216, ZN => n748);
   U903 : AOI221_X1 port map( B1 => n950, B2 => n221, C1 => n929, C2 => n223, A
                           => n951, ZN => n914);
   U904 : OAI222_X1 port map( A1 => n231, A2 => n905, B1 => n753, B2 => n228, 
                           C1 => n12, C2 => n952, ZN => n951);
   U905 : INV_X1 port map( A => n903, ZN => n753);
   U906 : OAI221_X1 port map( B1 => n953, B2 => n92, C1 => n932, C2 => n94, A 
                           => n954, ZN => n903);
   U907 : AOI222_X1 port map( A1 => n7, A2 => n955, B1 => n906, B2 => n375, C1 
                           => n376, C2 => n956, ZN => n954);
   U908 : INV_X1 port map( A => n756, ZN => n906);
   U909 : AOI222_X1 port map( A1 => n957, A2 => n16, B1 => n15, B2 => n920, C1 
                           => n936, C2 => n13, ZN => n756);
   U910 : OAI221_X1 port map( B1 => n165, B2 => n51, C1 => n52, C2 => n245, A 
                           => n958, ZN => n920);
   U911 : AOI222_X1 port map( A1 => DATA1(26), A2 => n17, B1 => DATA1(27), B2 
                           => n247, C1 => DATA1(23), C2 => n18, ZN => n958);
   U912 : INV_X1 port map( A => DATA1(25), ZN => n52);
   U913 : INV_X1 port map( A => n959, ZN => n214);
   U914 : OAI222_X1 port map( A1 => n219, A2 => n928, B1 => n949, B2 => n216, 
                           C1 => n960, C2 => n10, ZN => n891);
   U915 : AOI221_X1 port map( B1 => n961, B2 => n221, C1 => n950, C2 => n223, A
                           => n962, ZN => n928);
   U916 : OAI222_X1 port map( A1 => n231, A2 => n917, B1 => n905, B2 => n228, 
                           C1 => n12, C2 => n963, ZN => n962);
   U917 : INV_X1 port map( A => n915, ZN => n905);
   U918 : OAI221_X1 port map( B1 => n964, B2 => n92, C1 => n953, C2 => n94, A 
                           => n965, ZN => n915);
   U919 : AOI222_X1 port map( A1 => n7, A2 => n919, B1 => n375, B2 => n955, C1 
                           => n376, C2 => n966, ZN => n965);
   U920 : INV_X1 port map( A => n908, ZN => n955);
   U921 : AOI222_X1 port map( A1 => n15, A2 => n936, B1 => n967, B2 => n16, C1 
                           => n957, C2 => n13, ZN => n908);
   U922 : OAI221_X1 port map( B1 => n165, B2 => n50, C1 => n245, C2 => n51, A 
                           => n968, ZN => n936);
   U923 : AOI222_X1 port map( A1 => n17, A2 => DATA1(25), B1 => DATA1(26), B2 
                           => n247, C1 => DATA1(22), C2 => n18, ZN => n968);
   U924 : INV_X1 port map( A => DATA1(24), ZN => n51);
   U925 : INV_X1 port map( A => n670, ZN => n209);
   U926 : NAND2_X1 port map( A1 => n959, A2 => n969, ZN => n670);
   U927 : INV_X1 port map( A => n564, ZN => n207);
   U928 : NOR2_X1 port map( A1 => n970, A2 => n969, ZN => n564);
   U929 : OAI21_X1 port map( B1 => n925, B2 => n780, A => n959, ZN => n969);
   U930 : NOR2_X1 port map( A1 => n201, A2 => n860, ZN => n959);
   U931 : INV_X1 port map( A => n923, ZN => n201);
   U932 : NAND2_X1 port map( A1 => DATA2(3), A2 => n971, ZN => n923);
   U933 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(4), ZN => n780);
   U934 : INV_X1 port map( A => n878, ZN => n926);
   U935 : OAI222_X1 port map( A1 => n939, A2 => n10, B1 => n219, B2 => n949, C1
                           => n960, C2 => n216, ZN => n878);
   U936 : AOI221_X1 port map( B1 => n972, B2 => n221, C1 => n961, C2 => n223, A
                           => n973, ZN => n949);
   U937 : OAI222_X1 port map( A1 => n231, A2 => n931, B1 => n917, B2 => n228, 
                           C1 => n12, C2 => n942, ZN => n973);
   U938 : INV_X1 port map( A => n929, ZN => n917);
   U939 : OAI221_X1 port map( B1 => n974, B2 => n92, C1 => n964, C2 => n94, A 
                           => n975, ZN => n929);
   U940 : AOI222_X1 port map( A1 => n7, A2 => n934, B1 => n375, B2 => n919, C1 
                           => n376, C2 => n976, ZN => n975);
   U941 : INV_X1 port map( A => n932, ZN => n919);
   U942 : AOI222_X1 port map( A1 => n15, A2 => n957, B1 => n977, B2 => n16, C1 
                           => n967, C2 => n13, ZN => n932);
   U943 : OAI221_X1 port map( B1 => n165, B2 => n49, C1 => n245, C2 => n50, A 
                           => n978, ZN => n957);
   U944 : AOI222_X1 port map( A1 => DATA1(24), A2 => n17, B1 => DATA1(25), B2 
                           => n247, C1 => DATA1(21), C2 => n18, ZN => n978);
   U945 : INV_X1 port map( A => DATA1(23), ZN => n50);
   U946 : NAND2_X1 port map( A1 => n971, A2 => n979, ZN => n970);
   U947 : INV_X1 port map( A => n212, ZN => n617);
   U948 : NAND3_X1 port map( A1 => n980, A2 => n773, A3 => n925, ZN => n979);
   U949 : INV_X1 port map( A => n865, ZN => n889);
   U950 : OAI222_X1 port map( A1 => n219, A2 => n960, B1 => n939, B2 => n216, 
                           C1 => n892, C2 => n10, ZN => n865);
   U951 : AOI221_X1 port map( B1 => n940, B2 => n221, C1 => n981, C2 => n223, A
                           => n982, ZN => n892);
   U952 : OAI222_X1 port map( A1 => n231, A2 => n942, B1 => n228, B2 => n963, 
                           C1 => n12, C2 => n869, ZN => n982);
   U953 : INV_X1 port map( A => n893, ZN => n869);
   U954 : OAI221_X1 port map( B1 => n884, B2 => n92, C1 => n897, C2 => n94, A 
                           => n983, ZN => n893);
   U955 : AOI222_X1 port map( A1 => n7, A2 => n945, B1 => n375, B2 => n984, C1 
                           => n376, C2 => n871, ZN => n983);
   U956 : INV_X1 port map( A => n883, ZN => n871);
   U957 : AOI222_X1 port map( A1 => n15, A2 => n985, B1 => n898, B2 => n16, C1 
                           => n947, C2 => n13, ZN => n883);
   U958 : OAI221_X1 port map( B1 => n86, B2 => n165, C1 => n245, C2 => n676, A 
                           => n986, ZN => n898);
   U959 : AOI222_X1 port map( A1 => DATA1(11), A2 => n17, B1 => DATA1(12), B2 
                           => n247, C1 => DATA1(8), C2 => n18, ZN => n986);
   U960 : INV_X1 port map( A => DATA1(9), ZN => n86);
   U961 : INV_X1 port map( A => n987, ZN => n942);
   U962 : INV_X1 port map( A => n881, ZN => n940);
   U963 : OAI21_X1 port map( B1 => n764, B2 => n988, A => n219, ZN => n218);
   U964 : AOI221_X1 port map( B1 => n981, B2 => n221, C1 => n987, C2 => n223, A
                           => n989, ZN => n939);
   U965 : OAI222_X1 port map( A1 => n231, A2 => n963, B1 => n228, B2 => n952, 
                           C1 => n12, C2 => n881, ZN => n989);
   U966 : AOI221_X1 port map( B1 => n944, B2 => n68, C1 => n945, C2 => n70, A 
                           => n990, ZN => n881);
   U967 : OAI222_X1 port map( A1 => n2, A2 => n991, B1 => n237, B2 => n992, C1 
                           => n65, C2 => n884, ZN => n990);
   U968 : AOI222_X1 port map( A1 => n15, A2 => n993, B1 => n947, B2 => n16, C1 
                           => n985, C2 => n13, ZN => n884);
   U969 : OAI221_X1 port map( B1 => n165, B2 => n676, C1 => n245, C2 => n662, A
                           => n994, ZN => n947);
   U970 : AOI222_X1 port map( A1 => DATA1(12), A2 => n17, B1 => DATA1(13), B2 
                           => n247, C1 => DATA1(9), C2 => n18, ZN => n994);
   U971 : INV_X1 port map( A => DATA1(10), ZN => n676);
   U972 : INV_X1 port map( A => n375, ZN => n237);
   U973 : INV_X1 port map( A => n94, ZN => n70);
   U974 : INV_X1 port map( A => n92, ZN => n68);
   U975 : INV_X1 port map( A => n972, ZN => n963);
   U976 : AOI221_X1 port map( B1 => n987, B2 => n221, C1 => n972, C2 => n223, A
                           => n995, ZN => n960);
   U977 : OAI222_X1 port map( A1 => n231, A2 => n952, B1 => n228, B2 => n931, 
                           C1 => n12, C2 => n895, ZN => n995);
   U978 : INV_X1 port map( A => n981, ZN => n895);
   U979 : OAI221_X1 port map( B1 => n996, B2 => n92, C1 => n991, C2 => n94, A 
                           => n997, ZN => n981);
   U980 : AOI222_X1 port map( A1 => n7, A2 => n998, B1 => n375, B2 => n999, C1 
                           => n376, C2 => n944, ZN => n997);
   U981 : INV_X1 port map( A => n897, ZN => n944);
   U982 : AOI222_X1 port map( A1 => n15, A2 => n1000, B1 => n985, B2 => n16, C1
                           => n993, C2 => n13, ZN => n897);
   U983 : OAI221_X1 port map( B1 => n165, B2 => n662, C1 => n245, C2 => n641, A
                           => n1001, ZN => n985);
   U984 : AOI222_X1 port map( A1 => DATA1(13), A2 => n17, B1 => DATA1(14), B2 
                           => n247, C1 => DATA1(10), C2 => n18, ZN => n1001);
   U985 : INV_X1 port map( A => DATA1(11), ZN => n662);
   U986 : INV_X1 port map( A => n950, ZN => n931);
   U987 : OAI221_X1 port map( B1 => n1002, B2 => n92, C1 => n974, C2 => n94, A 
                           => n1003, ZN => n950);
   U988 : AOI222_X1 port map( A1 => n7, A2 => n956, B1 => n375, B2 => n934, C1 
                           => n376, C2 => n999, ZN => n1003);
   U989 : INV_X1 port map( A => n953, ZN => n934);
   U990 : AOI222_X1 port map( A1 => n15, A2 => n967, B1 => n1004, B2 => n16, C1
                           => n977, C2 => n13, ZN => n953);
   U991 : OAI221_X1 port map( B1 => n165, B2 => n48, C1 => n245, C2 => n49, A 
                           => n1005, ZN => n967);
   U992 : AOI222_X1 port map( A1 => DATA1(23), A2 => n17, B1 => DATA1(24), B2 
                           => n247, C1 => DATA1(20), C2 => n18, ZN => n1005);
   U993 : INV_X1 port map( A => DATA1(22), ZN => n49);
   U994 : INV_X1 port map( A => n961, ZN => n952);
   U995 : OAI221_X1 port map( B1 => n1006, B2 => n92, C1 => n1002, C2 => n94, A
                           => n1007, ZN => n961);
   U996 : AOI222_X1 port map( A1 => n7, A2 => n966, B1 => n375, B2 => n956, C1 
                           => n376, C2 => n998, ZN => n1007);
   U997 : INV_X1 port map( A => n992, ZN => n998);
   U998 : INV_X1 port map( A => n964, ZN => n956);
   U999 : AOI222_X1 port map( A1 => n15, A2 => n977, B1 => n1008, B2 => n16, C1
                           => n1004, C2 => n13, ZN => n964);
   U1000 : OAI221_X1 port map( B1 => n165, B2 => n47, C1 => n245, C2 => n48, A 
                           => n1009, ZN => n977);
   U1001 : AOI222_X1 port map( A1 => DATA1(22), A2 => n17, B1 => DATA1(23), B2 
                           => n247, C1 => DATA1(19), C2 => n18, ZN => n1009);
   U1002 : INV_X1 port map( A => DATA1(21), ZN => n48);
   U1003 : OAI21_X1 port map( B1 => n773, B2 => n988, A => n228, ZN => n1010);
   U1004 : OAI21_X1 port map( B1 => n980, B2 => n764, A => n219, ZN => n274);
   U1005 : OAI221_X1 port map( B1 => n992, B2 => n92, C1 => n1006, C2 => n94, A
                           => n1012, ZN => n972);
   U1006 : AOI222_X1 port map( A1 => n7, A2 => n976, B1 => n375, B2 => n966, C1
                           => n376, C2 => n984, ZN => n1012);
   U1007 : INV_X1 port map( A => n991, ZN => n984);
   U1008 : INV_X1 port map( A => n974, ZN => n966);
   U1009 : AOI222_X1 port map( A1 => n15, A2 => n1004, B1 => n1013, B2 => n16, 
                           C1 => n1008, C2 => n13, ZN => n974);
   U1010 : OAI221_X1 port map( B1 => n165, B2 => n46, C1 => n245, C2 => n47, A 
                           => n1014, ZN => n1004);
   U1011 : AOI222_X1 port map( A1 => DATA1(21), A2 => n17, B1 => DATA1(22), B2 
                           => n247, C1 => DATA1(18), C2 => n18, ZN => n1014);
   U1012 : INV_X1 port map( A => DATA1(20), ZN => n47);
   U1013 : NAND2_X1 port map( A1 => n12, A2 => n1011, ZN => n316);
   U1014 : OAI21_X1 port map( B1 => n724, B2 => n764, A => n1011, ZN => n227);
   U1015 : OAI221_X1 port map( B1 => n991, B2 => n92, C1 => n992, C2 => n94, A 
                           => n1015, ZN => n987);
   U1016 : AOI222_X1 port map( A1 => n7, A2 => n999, B1 => n375, B2 => n976, C1
                           => n376, C2 => n945, ZN => n1015);
   U1017 : INV_X1 port map( A => n996, ZN => n945);
   U1018 : AOI222_X1 port map( A1 => n15, A2 => n1016, B1 => n993, B2 => n16, 
                           C1 => n1000, C2 => n13, ZN => n996);
   U1019 : OAI221_X1 port map( B1 => n165, B2 => n641, C1 => n245, C2 => n628, 
                           A => n1017, ZN => n993);
   U1020 : AOI222_X1 port map( A1 => DATA1(14), A2 => n17, B1 => DATA1(15), B2 
                           => n247, C1 => DATA1(11), C2 => n18, ZN => n1017);
   U1021 : INV_X1 port map( A => DATA1(12), ZN => n641);
   U1022 : INV_X1 port map( A => n1002, ZN => n976);
   U1023 : AOI222_X1 port map( A1 => n15, A2 => n1008, B1 => n1018, B2 => n16, 
                           C1 => n1013, C2 => n13, ZN => n1002);
   U1024 : OAI221_X1 port map( B1 => n165, B2 => n45, C1 => n245, C2 => n46, A 
                           => n1019, ZN => n1008);
   U1025 : AOI222_X1 port map( A1 => DATA1(20), A2 => n17, B1 => DATA1(21), B2 
                           => n247, C1 => DATA1(17), C2 => n18, ZN => n1019);
   U1026 : INV_X1 port map( A => DATA1(19), ZN => n46);
   U1027 : INV_X1 port map( A => n1006, ZN => n999);
   U1028 : AOI222_X1 port map( A1 => n15, A2 => n1013, B1 => n1020, B2 => n16, 
                           C1 => n1018, C2 => n13, ZN => n1006);
   U1029 : OAI221_X1 port map( B1 => n165, B2 => n44, C1 => n245, C2 => n45, A 
                           => n1021, ZN => n1013);
   U1030 : AOI222_X1 port map( A1 => DATA1(19), A2 => n17, B1 => DATA1(20), B2 
                           => n247, C1 => DATA1(16), C2 => n18, ZN => n1021);
   U1031 : INV_X1 port map( A => DATA1(18), ZN => n45);
   U1032 : OAI21_X1 port map( B1 => DATA2(2), B2 => n971, A => n1023, ZN => 
                           n1011);
   U1033 : INV_X1 port map( A => n219, ZN => n971);
   U1034 : NAND2_X1 port map( A1 => n1023, A2 => n1024, ZN => n1022);
   U1035 : NAND4_X1 port map( A1 => n219, A2 => n724, A3 => n925, A4 => n980, 
                           ZN => n1024);
   U1036 : INV_X1 port map( A => DATA2(0), ZN => n724);
   U1037 : AOI222_X1 port map( A1 => n15, A2 => n1018, B1 => n1016, B2 => n16, 
                           C1 => n1020, C2 => n13, ZN => n992);
   U1038 : OAI221_X1 port map( B1 => n165, B2 => n43, C1 => n245, C2 => n44, A 
                           => n1025, ZN => n1018);
   U1039 : AOI222_X1 port map( A1 => DATA1(18), A2 => n17, B1 => DATA1(19), B2 
                           => n247, C1 => DATA1(15), C2 => n18, ZN => n1025);
   U1040 : INV_X1 port map( A => DATA1(17), ZN => n44);
   U1041 : INV_X1 port map( A => n376, ZN => n65);
   U1042 : AOI222_X1 port map( A1 => n15, A2 => n1020, B1 => n1000, B2 => n16, 
                           C1 => n1016, C2 => n13, ZN => n991);
   U1043 : OAI221_X1 port map( B1 => n165, B2 => n608, C1 => n245, C2 => n589, 
                           A => n1028, ZN => n1016);
   U1044 : AOI222_X1 port map( A1 => DATA1(16), A2 => n17, B1 => DATA1(17), B2 
                           => n247, C1 => DATA1(13), C2 => n18, ZN => n1028);
   U1045 : INV_X1 port map( A => n988, ZN => n1027);
   U1046 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(2), ZN => n988);
   U1047 : OAI221_X1 port map( B1 => n165, B2 => n628, C1 => n245, C2 => n608, 
                           A => n1029, ZN => n1000);
   U1048 : AOI222_X1 port map( A1 => DATA1(15), A2 => n17, B1 => DATA1(16), B2 
                           => n247, C1 => DATA1(12), C2 => n18, ZN => n1029);
   U1049 : INV_X1 port map( A => DATA1(14), ZN => n608);
   U1050 : INV_X1 port map( A => DATA1(13), ZN => n628);
   U1051 : OAI221_X1 port map( B1 => n165, B2 => n589, C1 => n245, C2 => n43, A
                           => n1030, ZN => n1020);
   U1052 : AOI222_X1 port map( A1 => DATA1(17), A2 => n17, B1 => DATA1(18), B2 
                           => n247, C1 => DATA1(14), C2 => n18, ZN => n1030);
   U1053 : INV_X1 port map( A => DATA1(16), ZN => n43);
   U1054 : AOI21_X1 port map( B1 => DATA2(1), B2 => DATA2(0), A => n247, ZN => 
                           n1031);
   U1055 : INV_X1 port map( A => DATA1(15), ZN => n589);
   U1056 : NOR2_X1 port map( A1 => n1032, A2 => n18, ZN => n534);
   U1057 : OR2_X1 port map( A1 => n247, A2 => DATA2(1), ZN => n1032);
   U1058 : OAI21_X1 port map( B1 => n925, B2 => n980, A => n1026, ZN => n242);
   U1059 : INV_X1 port map( A => n1023, ZN => n1026);
   U1060 : NAND2_X1 port map( A1 => n219, A2 => n773, ZN => n1023);
   U1061 : INV_X1 port map( A => DATA2(3), ZN => n773);
   U1062 : INV_X1 port map( A => DATA2(2), ZN => n980);
   U1063 : INV_X1 port map( A => DATA2(1), ZN => n925);
   U1064 : INV_X1 port map( A => n765, ZN => n1033);
   U1065 : NAND2_X1 port map( A1 => n860, A2 => DATA2(3), ZN => n765);
   U1066 : AND2_X1 port map( A1 => DATA2(4), A2 => DATA2(2), ZN => n860);
   U1067 : INV_X1 port map( A => n764, ZN => n859);
   U1068 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(1), ZN => n764);
   U1069 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(31), Z => N2548);
   U1070 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(30), Z => N2547);
   U1071 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(29), Z => N2546);
   U1072 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(28), Z => N2545);
   U1073 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(27), Z => N2544);
   U1074 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(26), Z => N2543);
   U1075 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(25), Z => N2542);
   U1076 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(24), Z => N2541);
   U1077 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(23), Z => N2540);
   U1078 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(22), Z => N2539);
   U1079 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(21), Z => N2538);
   U1080 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(20), Z => N2537);
   U1081 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(19), Z => N2536);
   U1082 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(18), Z => N2535);
   U1083 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(17), Z => N2534);
   U1084 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(16), Z => N2533);
   U1085 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(15), Z => N2532);
   U1086 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(14), Z => N2531);
   U1087 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(13), Z => N2530);
   U1088 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(12), Z => N2529);
   U1089 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(11), Z => N2528);
   U1090 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(10), Z => N2527);
   U1091 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(9), Z => N2526);
   U1092 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(8), Z => N2525);
   U1093 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(7), Z => N2524);
   U1094 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(6), Z => N2523);
   U1095 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(5), Z => N2522);
   U1096 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(4), Z => N2521);
   U1097 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(3), Z => N2520);
   U1098 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(2), Z => N2519);
   U1099 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(1), Z => N2518);
   U1100 : MUX2_X1 port map( A => n27, B => n28, S => DATA2(0), Z => N2517);
   U1101 : INV_X1 port map( A => FUNC(3), ZN => n723);
   U1102 : INV_X1 port map( A => FUNC(2), ZN => n726);
   U1103 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n728);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n1 is

   port( clk, reset, d : in std_logic;  Q : out std_logic);

end reg_nbit_n1;

architecture SYN_struc of reg_nbit_n1 is

   component FD_1911
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;

begin
   
   D_I_0 : FD_1911 port map( D => d, CK => clk, RESET => reset, Q => Q);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity check_branch_logic_N32 is

   port( input_val : in std_logic_vector (31 downto 0);  enable : in std_logic;
         decision : out std_logic);

end check_branch_logic_N32;

architecture SYN_behavioural of check_branch_logic_N32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U2 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => decision);
   U3 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U4 : NOR4_X1 port map( A1 => input_val(22), A2 => input_val(21), A3 => 
                           input_val(20), A4 => input_val(1), ZN => n6);
   U5 : NOR4_X1 port map( A1 => input_val(19), A2 => input_val(18), A3 => 
                           input_val(17), A4 => input_val(16), ZN => n5);
   U6 : NOR4_X1 port map( A1 => input_val(15), A2 => input_val(14), A3 => 
                           input_val(13), A4 => input_val(12), ZN => n4);
   U7 : NOR4_X1 port map( A1 => input_val(11), A2 => input_val(10), A3 => 
                           input_val(0), A4 => n7, ZN => n3);
   U8 : INV_X1 port map( A => enable, ZN => n7);
   U9 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n1);
   U10 : NOR4_X1 port map( A1 => n12, A2 => input_val(7), A3 => input_val(9), 
                           A4 => input_val(8), ZN => n11);
   U11 : OR2_X1 port map( A1 => input_val(6), A2 => input_val(5), ZN => n12);
   U12 : NOR4_X1 port map( A1 => input_val(4), A2 => input_val(3), A3 => 
                           input_val(31), A4 => input_val(30), ZN => n10);
   U13 : NOR4_X1 port map( A1 => input_val(2), A2 => input_val(29), A3 => 
                           input_val(28), A4 => input_val(27), ZN => n9);
   U14 : NOR4_X1 port map( A1 => input_val(26), A2 => input_val(25), A3 => 
                           input_val(24), A4 => input_val(23), ZN => n8);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n33_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (32 downto 0);  Q 
         : out std_logic_vector (32 downto 0));

end reg_nbit_n33_0;

architecture SYN_struc of reg_nbit_n33_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_1945
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1946
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1947
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1948
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1949
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1950
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1951
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1952
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1953
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1954
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1955
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1956
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1957
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1958
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1959
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1960
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1961
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1962
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1963
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1964
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1965
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1966
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1967
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1968
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1969
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1970
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1971
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1972
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1973
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1974
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1975
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1976
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_1977
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   D_I_0 : FD_1977 port map( D => d(0), CK => n4, RESET => n1, Q => Q(0));
   D_I_1 : FD_1976 port map( D => d(1), CK => n4, RESET => n1, Q => Q(1));
   D_I_2 : FD_1975 port map( D => d(2), CK => n4, RESET => n1, Q => Q(2));
   D_I_3 : FD_1974 port map( D => d(3), CK => n4, RESET => n1, Q => Q(3));
   D_I_4 : FD_1973 port map( D => d(4), CK => n4, RESET => n1, Q => Q(4));
   D_I_5 : FD_1972 port map( D => d(5), CK => n4, RESET => n1, Q => Q(5));
   D_I_6 : FD_1971 port map( D => d(6), CK => n4, RESET => n1, Q => Q(6));
   D_I_7 : FD_1970 port map( D => d(7), CK => n4, RESET => n1, Q => Q(7));
   D_I_8 : FD_1969 port map( D => d(8), CK => n4, RESET => n1, Q => Q(8));
   D_I_9 : FD_1968 port map( D => d(9), CK => n4, RESET => n1, Q => Q(9));
   D_I_10 : FD_1967 port map( D => d(10), CK => n4, RESET => n1, Q => Q(10));
   D_I_11 : FD_1966 port map( D => d(11), CK => n5, RESET => n1, Q => Q(11));
   D_I_12 : FD_1965 port map( D => d(12), CK => n5, RESET => n2, Q => Q(12));
   D_I_13 : FD_1964 port map( D => d(13), CK => n5, RESET => n2, Q => Q(13));
   D_I_14 : FD_1963 port map( D => d(14), CK => n5, RESET => n2, Q => Q(14));
   D_I_15 : FD_1962 port map( D => d(15), CK => n5, RESET => n2, Q => Q(15));
   D_I_16 : FD_1961 port map( D => d(16), CK => n5, RESET => n2, Q => Q(16));
   D_I_17 : FD_1960 port map( D => d(17), CK => n5, RESET => n2, Q => Q(17));
   D_I_18 : FD_1959 port map( D => d(18), CK => n5, RESET => n2, Q => Q(18));
   D_I_19 : FD_1958 port map( D => d(19), CK => n5, RESET => n2, Q => Q(19));
   D_I_20 : FD_1957 port map( D => d(20), CK => n5, RESET => n2, Q => Q(20));
   D_I_21 : FD_1956 port map( D => d(21), CK => n5, RESET => n2, Q => Q(21));
   D_I_22 : FD_1955 port map( D => d(22), CK => n6, RESET => n2, Q => Q(22));
   D_I_23 : FD_1954 port map( D => d(23), CK => n6, RESET => n2, Q => Q(23));
   D_I_24 : FD_1953 port map( D => d(24), CK => n6, RESET => n3, Q => Q(24));
   D_I_25 : FD_1952 port map( D => d(25), CK => n6, RESET => n3, Q => Q(25));
   D_I_26 : FD_1951 port map( D => d(26), CK => n6, RESET => n3, Q => Q(26));
   D_I_27 : FD_1950 port map( D => d(27), CK => n6, RESET => n3, Q => Q(27));
   D_I_28 : FD_1949 port map( D => d(28), CK => n6, RESET => n3, Q => Q(28));
   D_I_29 : FD_1948 port map( D => d(29), CK => n6, RESET => n3, Q => Q(29));
   D_I_30 : FD_1947 port map( D => d(30), CK => n6, RESET => n3, Q => Q(30));
   D_I_31 : FD_1946 port map( D => d(31), CK => n6, RESET => n3, Q => Q(31));
   D_I_32 : FD_1945 port map( D => d(32), CK => n6, RESET => n3, Q => Q(32));
   U1 : BUF_X1 port map( A => reset, Z => n1);
   U2 : BUF_X1 port map( A => reset, Z => n2);
   U3 : BUF_X1 port map( A => reset, Z => n3);
   U4 : BUF_X1 port map( A => clk, Z => n4);
   U5 : BUF_X1 port map( A => clk, Z => n5);
   U6 : BUF_X1 port map( A => clk, Z => n6);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_zbit_nbit_N32_Z1_0 is

   port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_zbit_nbit_N32_Z1_0;

architecture SYN_beh of MUX_zbit_nbit_N32_Z1_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n34, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15
      , n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32 : std_logic;

begin
   
   Y_reg_31_inst : DLH_X1 port map( G => n34, D => n7, Q => Y(31));
   Y_reg_30_inst : DLH_X1 port map( G => n34, D => n8, Q => Y(30));
   Y_reg_29_inst : DLH_X1 port map( G => n34, D => n9, Q => Y(29));
   Y_reg_28_inst : DLH_X1 port map( G => n34, D => n10, Q => Y(28));
   Y_reg_27_inst : DLH_X1 port map( G => n34, D => n11, Q => Y(27));
   Y_reg_26_inst : DLH_X1 port map( G => n34, D => n13, Q => Y(26));
   Y_reg_25_inst : DLH_X1 port map( G => n34, D => n14, Q => Y(25));
   Y_reg_24_inst : DLH_X1 port map( G => n34, D => n15, Q => Y(24));
   Y_reg_23_inst : DLH_X1 port map( G => n34, D => n16, Q => Y(23));
   Y_reg_22_inst : DLH_X1 port map( G => n34, D => n17, Q => Y(22));
   Y_reg_21_inst : DLH_X1 port map( G => n34, D => n18, Q => Y(21));
   Y_reg_20_inst : DLH_X1 port map( G => n34, D => n19, Q => Y(20));
   Y_reg_19_inst : DLH_X1 port map( G => n34, D => n20, Q => Y(19));
   Y_reg_18_inst : DLH_X1 port map( G => n34, D => n21, Q => Y(18));
   Y_reg_17_inst : DLH_X1 port map( G => n34, D => n22, Q => Y(17));
   Y_reg_16_inst : DLH_X1 port map( G => n34, D => n23, Q => Y(16));
   Y_reg_15_inst : DLH_X1 port map( G => n34, D => n24, Q => Y(15));
   Y_reg_14_inst : DLH_X1 port map( G => n34, D => n25, Q => Y(14));
   Y_reg_13_inst : DLH_X1 port map( G => n34, D => n26, Q => Y(13));
   Y_reg_12_inst : DLH_X1 port map( G => n34, D => n27, Q => Y(12));
   Y_reg_11_inst : DLH_X1 port map( G => n34, D => n28, Q => Y(11));
   Y_reg_10_inst : DLH_X1 port map( G => n34, D => n29, Q => Y(10));
   Y_reg_9_inst : DLH_X1 port map( G => n34, D => n30, Q => Y(9));
   Y_reg_8_inst : DLH_X1 port map( G => n34, D => n31, Q => Y(8));
   Y_reg_7_inst : DLH_X1 port map( G => n34, D => n32, Q => Y(7));
   Y_reg_6_inst : DLH_X1 port map( G => n34, D => n1, Q => Y(6));
   Y_reg_5_inst : DLH_X1 port map( G => n34, D => n2, Q => Y(5));
   Y_reg_4_inst : DLH_X1 port map( G => n34, D => n3, Q => Y(4));
   Y_reg_3_inst : DLH_X1 port map( G => n34, D => n4, Q => Y(3));
   Y_reg_2_inst : DLH_X1 port map( G => n34, D => n5, Q => Y(2));
   Y_reg_1_inst : DLH_X1 port map( G => n34, D => n6, Q => Y(1));
   Y_reg_0_inst : DLH_X1 port map( G => n34, D => n12, Q => Y(0));
   n34 <= '1';
   U3 : MUX2_X1 port map( A => inputs(25), B => inputs(57), S => SEL, Z => n1);
   U4 : MUX2_X1 port map( A => inputs(26), B => inputs(58), S => SEL, Z => n2);
   U5 : MUX2_X1 port map( A => inputs(27), B => inputs(59), S => SEL, Z => n3);
   U6 : MUX2_X1 port map( A => inputs(28), B => inputs(60), S => SEL, Z => n4);
   U7 : MUX2_X1 port map( A => inputs(29), B => inputs(61), S => SEL, Z => n5);
   U8 : MUX2_X1 port map( A => inputs(30), B => inputs(62), S => SEL, Z => n6);
   U9 : MUX2_X1 port map( A => inputs(0), B => inputs(32), S => SEL, Z => n7);
   U10 : MUX2_X1 port map( A => inputs(1), B => inputs(33), S => SEL, Z => n8);
   U11 : MUX2_X1 port map( A => inputs(2), B => inputs(34), S => SEL, Z => n9);
   U12 : MUX2_X1 port map( A => inputs(3), B => inputs(35), S => SEL, Z => n10)
                           ;
   U13 : MUX2_X1 port map( A => inputs(4), B => inputs(36), S => SEL, Z => n11)
                           ;
   U14 : MUX2_X1 port map( A => inputs(31), B => inputs(63), S => SEL, Z => n12
                           );
   U15 : MUX2_X1 port map( A => inputs(5), B => inputs(37), S => SEL, Z => n13)
                           ;
   U16 : MUX2_X1 port map( A => inputs(6), B => inputs(38), S => SEL, Z => n14)
                           ;
   U17 : MUX2_X1 port map( A => inputs(7), B => inputs(39), S => SEL, Z => n15)
                           ;
   U18 : MUX2_X1 port map( A => inputs(8), B => inputs(40), S => SEL, Z => n16)
                           ;
   U19 : MUX2_X1 port map( A => inputs(9), B => inputs(41), S => SEL, Z => n17)
                           ;
   U20 : MUX2_X1 port map( A => inputs(10), B => inputs(42), S => SEL, Z => n18
                           );
   U21 : MUX2_X1 port map( A => inputs(11), B => inputs(43), S => SEL, Z => n19
                           );
   U22 : MUX2_X1 port map( A => inputs(12), B => inputs(44), S => SEL, Z => n20
                           );
   U23 : MUX2_X1 port map( A => inputs(13), B => inputs(45), S => SEL, Z => n21
                           );
   U24 : MUX2_X1 port map( A => inputs(14), B => inputs(46), S => SEL, Z => n22
                           );
   U25 : MUX2_X1 port map( A => inputs(15), B => inputs(47), S => SEL, Z => n23
                           );
   U26 : MUX2_X1 port map( A => inputs(16), B => inputs(48), S => SEL, Z => n24
                           );
   U27 : MUX2_X1 port map( A => inputs(17), B => inputs(49), S => SEL, Z => n25
                           );
   U28 : MUX2_X1 port map( A => inputs(18), B => inputs(50), S => SEL, Z => n26
                           );
   U29 : MUX2_X1 port map( A => inputs(19), B => inputs(51), S => SEL, Z => n27
                           );
   U30 : MUX2_X1 port map( A => inputs(20), B => inputs(52), S => SEL, Z => n28
                           );
   U31 : MUX2_X1 port map( A => inputs(21), B => inputs(53), S => SEL, Z => n29
                           );
   U32 : MUX2_X1 port map( A => inputs(22), B => inputs(54), S => SEL, Z => n30
                           );
   U33 : MUX2_X1 port map( A => inputs(23), B => inputs(55), S => SEL, Z => n31
                           );
   U34 : MUX2_X1 port map( A => inputs(24), B => inputs(56), S => SEL, Z => n32
                           );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_extension_N32_STARTING_BIT26 is

   port( val_to_exetend : in std_logic_vector (25 downto 0);  enable : in 
         std_logic;  extended_val : out std_logic_vector (31 downto 0));

end sign_extension_N32_STARTING_BIT26;

architecture SYN_behavioural of sign_extension_N32_STARTING_BIT26 is

   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;

begin
   
   extended_val_reg_31_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(31));
   extended_val_reg_30_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(30));
   extended_val_reg_29_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(29));
   extended_val_reg_28_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(28));
   extended_val_reg_27_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(27));
   extended_val_reg_26_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(26));
   extended_val_reg_25_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(25), Q => extended_val(25));
   extended_val_reg_24_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(24), Q => extended_val(24));
   extended_val_reg_23_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(23), Q => extended_val(23));
   extended_val_reg_22_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(22), Q => extended_val(22));
   extended_val_reg_21_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(21), Q => extended_val(21));
   extended_val_reg_20_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(20), Q => extended_val(20));
   extended_val_reg_19_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(19), Q => extended_val(19));
   extended_val_reg_18_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(18), Q => extended_val(18));
   extended_val_reg_17_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(17), Q => extended_val(17));
   extended_val_reg_16_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(16), Q => extended_val(16));
   extended_val_reg_15_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(15));
   extended_val_reg_14_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(14), Q => extended_val(14));
   extended_val_reg_13_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(13), Q => extended_val(13));
   extended_val_reg_12_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(12), Q => extended_val(12));
   extended_val_reg_11_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(11), Q => extended_val(11));
   extended_val_reg_10_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(10), Q => extended_val(10));
   extended_val_reg_9_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(9), Q => extended_val(9));
   extended_val_reg_8_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(8), Q => extended_val(8));
   extended_val_reg_7_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(7), Q => extended_val(7));
   extended_val_reg_6_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(6), Q => extended_val(6));
   extended_val_reg_5_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(5), Q => extended_val(5));
   extended_val_reg_4_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(4), Q => extended_val(4));
   extended_val_reg_3_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(3), Q => extended_val(3));
   extended_val_reg_2_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(2), Q => extended_val(2));
   extended_val_reg_1_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(1), Q => extended_val(1));
   extended_val_reg_0_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(0), Q => extended_val(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_extension_N32_STARTING_BIT16 is

   port( val_to_exetend : in std_logic_vector (15 downto 0);  enable : in 
         std_logic;  extended_val : out std_logic_vector (31 downto 0));

end sign_extension_N32_STARTING_BIT16;

architecture SYN_behavioural of sign_extension_N32_STARTING_BIT16 is

   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;

begin
   
   extended_val_reg_31_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(31));
   extended_val_reg_30_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(30));
   extended_val_reg_29_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(29));
   extended_val_reg_28_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(28));
   extended_val_reg_27_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(27));
   extended_val_reg_26_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(26));
   extended_val_reg_25_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(25));
   extended_val_reg_24_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(24));
   extended_val_reg_23_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(23));
   extended_val_reg_22_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(22));
   extended_val_reg_21_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(21));
   extended_val_reg_20_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(20));
   extended_val_reg_19_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(19));
   extended_val_reg_18_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(18));
   extended_val_reg_17_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(17));
   extended_val_reg_16_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(16));
   extended_val_reg_15_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(15), Q => extended_val(15));
   extended_val_reg_14_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(14), Q => extended_val(14));
   extended_val_reg_13_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(13), Q => extended_val(13));
   extended_val_reg_12_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(12), Q => extended_val(12));
   extended_val_reg_11_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(11), Q => extended_val(11));
   extended_val_reg_10_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(10), Q => extended_val(10));
   extended_val_reg_9_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(9), Q => extended_val(9));
   extended_val_reg_8_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(8), Q => extended_val(8));
   extended_val_reg_7_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(7), Q => extended_val(7));
   extended_val_reg_6_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(6), Q => extended_val(6));
   extended_val_reg_5_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(5), Q => extended_val(5));
   extended_val_reg_4_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(4), Q => extended_val(4));
   extended_val_reg_3_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(3), Q => extended_val(3));
   extended_val_reg_2_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(2), Q => extended_val(2));
   extended_val_reg_1_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(1), Q => extended_val(1));
   extended_val_reg_0_inst : DLH_X1 port map( G => enable, D => 
                           val_to_exetend(0), Q => extended_val(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, 
      N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55
      , N56, N57, N58, N59, N60, N61, N62, N96, N97, N98, N99, N100, N101, N102
      , N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
      N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, 
      N127, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, 
      N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, 
      N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, 
      N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, 
      N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, 
      N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, n1147, n1148, 
      n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
      n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
      n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
      n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
      n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, 
      n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31_port, n32_port, 
      n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, 
      n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, 
      n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, 
      n54_port, n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, 
      n61_port, n62_port, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73
      , n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, 
      n88, n89, n90, n91, n92, n93, n94, n95, n96_port, n97_port, n98_port, 
      n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114_port, n115_port, n116_port, 
      n117_port, n118_port, n119_port, n120_port, n121_port, n122_port, 
      n123_port, n124_port, n125_port, n126_port, n127_port, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385_port, n386_port, n387_port, n388_port, n389_port, 
      n390_port, n391_port, n392_port, n393_port, n394_port, n395_port, 
      n396_port, n397_port, n398_port, n399_port, n400_port, n401_port, 
      n402_port, n403_port, n404_port, n405_port, n406_port, n407_port, 
      n408_port, n409_port, n410_port, n411_port, n412_port, n413_port, 
      n414_port, n415_port, n416_port, n417_port, n418_port, n419_port, 
      n420_port, n421_port, n422_port, n423_port, n424_port, n425_port, 
      n426_port, n427_port, n428_port, n429_port, n430_port, n431_port, 
      n432_port, n433_port, n434_port, n435_port, n436_port, n437_port, 
      n438_port, n439_port, n440_port, n441_port, n442_port, n443_port, 
      n444_port, n445_port, n446_port, n447_port, n448_port, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n_4445, n_4446, 
      n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, 
      n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, 
      n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, 
      n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, 
      n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, 
      n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, 
      n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, 
      n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, 
      n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, 
      n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, 
      n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, 
      n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, 
      n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, 
      n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, 
      n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, 
      n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, 
      n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, 
      n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, 
      n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, 
      n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, 
      n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, 
      n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, 
      n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, 
      n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, 
      n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, 
      n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, 
      n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, 
      n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, 
      n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, 
      n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, 
      n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, 
      n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, 
      n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, 
      n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, 
      n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, 
      n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, 
      n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, 
      n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, 
      n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, 
      n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, 
      n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, 
      n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, 
      n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, 
      n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, 
      n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, 
      n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, 
      n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, 
      n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, 
      n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, 
      n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, 
      n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, 
      n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, 
      n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, 
      n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, 
      n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, 
      n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, 
      n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, 
      n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, 
      n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, 
      n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, 
      n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, 
      n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, 
      n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, 
      n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, 
      n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, 
      n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, 
      n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, 
      n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, 
      n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, 
      n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, 
      n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, 
      n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, 
      n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, 
      n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112, 
      n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, 
      n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, 
      n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, 
      n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, 
      n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5157, 
      n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, 
      n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, 
      n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, 
      n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, 
      n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, 
      n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, 
      n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220, 
      n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, 
      n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, 
      n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, 
      n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, 
      n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, 
      n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, 
      n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, 
      n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, 
      n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, 
      n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, 
      n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, 
      n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328, 
      n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337, 
      n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, 
      n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, 
      n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, 
      n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, 
      n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, 
      n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, 
      n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, 
      n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409, 
      n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416, n_5417, n_5418, 
      n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, 
      n_5428, n_5429, n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, 
      n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, 
      n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, 
      n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, 
      n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, 
      n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481, 
      n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489, n_5490, 
      n_5491, n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, 
      n_5500, n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, 
      n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, 
      n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, 
      n_5527, n_5528, n_5529, n_5530, n_5531, n_5532 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => n370, Q => 
                           REGISTERS_0_31_port, QN => n_4445);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => n373, Q => 
                           REGISTERS_0_30_port, QN => n_4446);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => n376, Q => 
                           REGISTERS_0_29_port, QN => n_4447);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => n379, Q => 
                           REGISTERS_0_28_port, QN => n_4448);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => n383, Q => 
                           REGISTERS_0_27_port, QN => n_4449);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => n364, Q => 
                           REGISTERS_0_26_port, QN => n_4450);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => n352, Q => 
                           REGISTERS_0_25_port, QN => n_4451);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => n355, Q => 
                           REGISTERS_0_24_port, QN => n_4452);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => n343, Q => 
                           REGISTERS_0_23_port, QN => n_4453);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => n346, Q => 
                           REGISTERS_0_22_port, QN => n_4454);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => n349, Q => 
                           REGISTERS_0_21_port, QN => n_4455);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => n330, Q => 
                           REGISTERS_0_20_port, QN => n_4456);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => n333, Q => 
                           REGISTERS_0_19_port, QN => n_4457);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => n336, Q => 
                           REGISTERS_0_18_port, QN => n_4458);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => n358, Q => 
                           REGISTERS_0_17_port, QN => n_4459);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => n340, Q => 
                           REGISTERS_0_16_port, QN => n_4460);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => n324, Q => 
                           REGISTERS_0_15_port, QN => n_4461);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => n327, Q => 
                           REGISTERS_0_14_port, QN => n_4462);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => n321, Q => 
                           REGISTERS_0_13_port, QN => n_4463);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => n318, Q => 
                           REGISTERS_0_12_port, QN => n_4464);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => n315, Q => 
                           REGISTERS_0_11_port, QN => n_4465);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => n312, Q => 
                           REGISTERS_0_10_port, QN => n_4466);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => n309, Q => 
                           REGISTERS_0_9_port, QN => n_4467);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => n306, Q => 
                           REGISTERS_0_8_port, QN => n_4468);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => n303, Q => 
                           REGISTERS_0_7_port, QN => n_4469);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => n299, Q => 
                           REGISTERS_0_6_port, QN => n_4470);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => n296, Q => 
                           REGISTERS_0_5_port, QN => n_4471);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => n293, Q => 
                           REGISTERS_0_4_port, QN => n_4472);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => n290, Q => 
                           REGISTERS_0_3_port, QN => n_4473);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => n361, Q => 
                           REGISTERS_0_2_port, QN => n_4474);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => n287, Q => 
                           REGISTERS_0_1_port, QN => n_4475);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => n367, Q => 
                           REGISTERS_0_0_port, QN => n_4476);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => n370, Q => 
                           REGISTERS_1_31_port, QN => n_4477);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => n373, Q => 
                           REGISTERS_1_30_port, QN => n_4478);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => n376, Q => 
                           REGISTERS_1_29_port, QN => n_4479);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => n380, Q => 
                           REGISTERS_1_28_port, QN => n_4480);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => n383, Q => 
                           REGISTERS_1_27_port, QN => n_4481);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => n364, Q => 
                           REGISTERS_1_26_port, QN => n_4482);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => n352, Q => 
                           REGISTERS_1_25_port, QN => n_4483);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => n355, Q => 
                           REGISTERS_1_24_port, QN => n_4484);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => n343, Q => 
                           REGISTERS_1_23_port, QN => n_4485);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => n346, Q => 
                           REGISTERS_1_22_port, QN => n_4486);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => n349, Q => 
                           REGISTERS_1_21_port, QN => n_4487);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => n330, Q => 
                           REGISTERS_1_20_port, QN => n_4488);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => n333, Q => 
                           REGISTERS_1_19_port, QN => n_4489);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => n337, Q => 
                           REGISTERS_1_18_port, QN => n_4490);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => n358, Q => 
                           REGISTERS_1_17_port, QN => n_4491);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => n340, Q => 
                           REGISTERS_1_16_port, QN => n_4492);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => n324, Q => 
                           REGISTERS_1_15_port, QN => n_4493);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => n327, Q => 
                           REGISTERS_1_14_port, QN => n_4494);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => n321, Q => 
                           REGISTERS_1_13_port, QN => n_4495);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => n318, Q => 
                           REGISTERS_1_12_port, QN => n_4496);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => n315, Q => 
                           REGISTERS_1_11_port, QN => n_4497);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => n312, Q => 
                           REGISTERS_1_10_port, QN => n_4498);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => n309, Q => 
                           REGISTERS_1_9_port, QN => n_4499);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => n306, Q => 
                           REGISTERS_1_8_port, QN => n_4500);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => n303, Q => 
                           REGISTERS_1_7_port, QN => n_4501);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => n300, Q => 
                           REGISTERS_1_6_port, QN => n_4502);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => n296, Q => 
                           REGISTERS_1_5_port, QN => n_4503);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => n293, Q => 
                           REGISTERS_1_4_port, QN => n_4504);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => n290, Q => 
                           REGISTERS_1_3_port, QN => n_4505);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => n361, Q => 
                           REGISTERS_1_2_port, QN => n_4506);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => n287, Q => 
                           REGISTERS_1_1_port, QN => n_4507);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => n367, Q => 
                           REGISTERS_1_0_port, QN => n_4508);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => n370, Q => 
                           REGISTERS_2_31_port, QN => n_4509);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => n373, Q => 
                           REGISTERS_2_30_port, QN => n_4510);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => n377, Q => 
                           REGISTERS_2_29_port, QN => n_4511);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => n380, Q => 
                           REGISTERS_2_28_port, QN => n_4512);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => n383, Q => 
                           REGISTERS_2_27_port, QN => n_4513);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => n364, Q => 
                           REGISTERS_2_26_port, QN => n_4514);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => n352, Q => 
                           REGISTERS_2_25_port, QN => n_4515);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => n355, Q => 
                           REGISTERS_2_24_port, QN => n_4516);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => n343, Q => 
                           REGISTERS_2_23_port, QN => n_4517);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => n346, Q => 
                           REGISTERS_2_22_port, QN => n_4518);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => n349, Q => 
                           REGISTERS_2_21_port, QN => n_4519);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => n330, Q => 
                           REGISTERS_2_20_port, QN => n_4520);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => n334, Q => 
                           REGISTERS_2_19_port, QN => n_4521);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => n337, Q => 
                           REGISTERS_2_18_port, QN => n_4522);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => n358, Q => 
                           REGISTERS_2_17_port, QN => n_4523);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => n340, Q => 
                           REGISTERS_2_16_port, QN => n_4524);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => n324, Q => 
                           REGISTERS_2_15_port, QN => n_4525);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => n327, Q => 
                           REGISTERS_2_14_port, QN => n_4526);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => n321, Q => 
                           REGISTERS_2_13_port, QN => n_4527);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => n318, Q => 
                           REGISTERS_2_12_port, QN => n_4528);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => n315, Q => 
                           REGISTERS_2_11_port, QN => n_4529);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => n312, Q => 
                           REGISTERS_2_10_port, QN => n_4530);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => n309, Q => 
                           REGISTERS_2_9_port, QN => n_4531);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => n306, Q => 
                           REGISTERS_2_8_port, QN => n_4532);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => n303, Q => 
                           REGISTERS_2_7_port, QN => n_4533);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => n300, Q => 
                           REGISTERS_2_6_port, QN => n_4534);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => n297, Q => 
                           REGISTERS_2_5_port, QN => n_4535);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => n293, Q => 
                           REGISTERS_2_4_port, QN => n_4536);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => n290, Q => 
                           REGISTERS_2_3_port, QN => n_4537);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => n361, Q => 
                           REGISTERS_2_2_port, QN => n_4538);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => n287, Q => 
                           REGISTERS_2_1_port, QN => n_4539);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => n367, Q => 
                           REGISTERS_2_0_port, QN => n_4540);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => n370, Q => 
                           REGISTERS_3_31_port, QN => n_4541);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => n374, Q => 
                           REGISTERS_3_30_port, QN => n_4542);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => n377, Q => 
                           REGISTERS_3_29_port, QN => n_4543);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => n380, Q => 
                           REGISTERS_3_28_port, QN => n_4544);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => n383, Q => 
                           REGISTERS_3_27_port, QN => n_4545);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => n364, Q => 
                           REGISTERS_3_26_port, QN => n_4546);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => n352, Q => 
                           REGISTERS_3_25_port, QN => n_4547);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => n355, Q => 
                           REGISTERS_3_24_port, QN => n_4548);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => n343, Q => 
                           REGISTERS_3_23_port, QN => n_4549);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => n346, Q => 
                           REGISTERS_3_22_port, QN => n_4550);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => n349, Q => 
                           REGISTERS_3_21_port, QN => n_4551);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => n331, Q => 
                           REGISTERS_3_20_port, QN => n_4552);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => n334, Q => 
                           REGISTERS_3_19_port, QN => n_4553);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => n337, Q => 
                           REGISTERS_3_18_port, QN => n_4554);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => n358, Q => 
                           REGISTERS_3_17_port, QN => n_4555);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => n340, Q => 
                           REGISTERS_3_16_port, QN => n_4556);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => n324, Q => 
                           REGISTERS_3_15_port, QN => n_4557);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => n328, Q => 
                           REGISTERS_3_14_port, QN => n_4558);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => n321, Q => 
                           REGISTERS_3_13_port, QN => n_4559);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => n318, Q => 
                           REGISTERS_3_12_port, QN => n_4560);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => n315, Q => 
                           REGISTERS_3_11_port, QN => n_4561);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => n312, Q => 
                           REGISTERS_3_10_port, QN => n_4562);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => n309, Q => 
                           REGISTERS_3_9_port, QN => n_4563);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => n306, Q => 
                           REGISTERS_3_8_port, QN => n_4564);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => n303, Q => 
                           REGISTERS_3_7_port, QN => n_4565);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => n300, Q => 
                           REGISTERS_3_6_port, QN => n_4566);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => n297, Q => 
                           REGISTERS_3_5_port, QN => n_4567);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => n294, Q => 
                           REGISTERS_3_4_port, QN => n_4568);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => n290, Q => 
                           REGISTERS_3_3_port, QN => n_4569);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => n361, Q => 
                           REGISTERS_3_2_port, QN => n_4570);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => n287, Q => 
                           REGISTERS_3_1_port, QN => n_4571);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => n367, Q => 
                           REGISTERS_3_0_port, QN => n_4572);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => n371, Q => 
                           REGISTERS_4_31_port, QN => n_4573);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => n374, Q => 
                           REGISTERS_4_30_port, QN => n_4574);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => n377, Q => 
                           REGISTERS_4_29_port, QN => n_4575);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => n380, Q => 
                           REGISTERS_4_28_port, QN => n_4576);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => n383, Q => 
                           REGISTERS_4_27_port, QN => n_4577);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => n364, Q => 
                           REGISTERS_4_26_port, QN => n_4578);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => n352, Q => 
                           REGISTERS_4_25_port, QN => n_4579);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => n355, Q => 
                           REGISTERS_4_24_port, QN => n_4580);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => n343, Q => 
                           REGISTERS_4_23_port, QN => n_4581);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => n346, Q => 
                           REGISTERS_4_22_port, QN => n_4582);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => n349, Q => 
                           REGISTERS_4_21_port, QN => n_4583);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => n331, Q => 
                           REGISTERS_4_20_port, QN => n_4584);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => n334, Q => 
                           REGISTERS_4_19_port, QN => n_4585);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => n337, Q => 
                           REGISTERS_4_18_port, QN => n_4586);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => n358, Q => 
                           REGISTERS_4_17_port, QN => n_4587);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => n340, Q => 
                           REGISTERS_4_16_port, QN => n_4588);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => n325, Q => 
                           REGISTERS_4_15_port, QN => n_4589);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => n328, Q => 
                           REGISTERS_4_14_port, QN => n_4590);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => n321, Q => 
                           REGISTERS_4_13_port, QN => n_4591);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => n318, Q => 
                           REGISTERS_4_12_port, QN => n_4592);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => n315, Q => 
                           REGISTERS_4_11_port, QN => n_4593);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => n312, Q => 
                           REGISTERS_4_10_port, QN => n_4594);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => n309, Q => 
                           REGISTERS_4_9_port, QN => n_4595);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => n306, Q => 
                           REGISTERS_4_8_port, QN => n_4596);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => n303, Q => 
                           REGISTERS_4_7_port, QN => n_4597);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => n300, Q => 
                           REGISTERS_4_6_port, QN => n_4598);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => n297, Q => 
                           REGISTERS_4_5_port, QN => n_4599);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => n294, Q => 
                           REGISTERS_4_4_port, QN => n_4600);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => n291, Q => 
                           REGISTERS_4_3_port, QN => n_4601);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => n361, Q => 
                           REGISTERS_4_2_port, QN => n_4602);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => n287, Q => 
                           REGISTERS_4_1_port, QN => n_4603);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => n367, Q => 
                           REGISTERS_4_0_port, QN => n_4604);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => n371, Q => 
                           REGISTERS_5_31_port, QN => n_4605);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => n374, Q => 
                           REGISTERS_5_30_port, QN => n_4606);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => n377, Q => 
                           REGISTERS_5_29_port, QN => n_4607);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => n380, Q => 
                           REGISTERS_5_28_port, QN => n_4608);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => n383, Q => 
                           REGISTERS_5_27_port, QN => n_4609);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => n364, Q => 
                           REGISTERS_5_26_port, QN => n_4610);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => n352, Q => 
                           REGISTERS_5_25_port, QN => n_4611);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => n355, Q => 
                           REGISTERS_5_24_port, QN => n_4612);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => n343, Q => 
                           REGISTERS_5_23_port, QN => n_4613);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => n346, Q => 
                           REGISTERS_5_22_port, QN => n_4614);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => n349, Q => 
                           REGISTERS_5_21_port, QN => n_4615);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => n331, Q => 
                           REGISTERS_5_20_port, QN => n_4616);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => n334, Q => 
                           REGISTERS_5_19_port, QN => n_4617);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => n337, Q => 
                           REGISTERS_5_18_port, QN => n_4618);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => n358, Q => 
                           REGISTERS_5_17_port, QN => n_4619);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => n340, Q => 
                           REGISTERS_5_16_port, QN => n_4620);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => n325, Q => 
                           REGISTERS_5_15_port, QN => n_4621);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => n328, Q => 
                           REGISTERS_5_14_port, QN => n_4622);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => n322, Q => 
                           REGISTERS_5_13_port, QN => n_4623);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => n318, Q => 
                           REGISTERS_5_12_port, QN => n_4624);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => n315, Q => 
                           REGISTERS_5_11_port, QN => n_4625);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => n312, Q => 
                           REGISTERS_5_10_port, QN => n_4626);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => n309, Q => 
                           REGISTERS_5_9_port, QN => n_4627);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => n306, Q => 
                           REGISTERS_5_8_port, QN => n_4628);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => n303, Q => 
                           REGISTERS_5_7_port, QN => n_4629);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => n300, Q => 
                           REGISTERS_5_6_port, QN => n_4630);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => n297, Q => 
                           REGISTERS_5_5_port, QN => n_4631);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => n294, Q => 
                           REGISTERS_5_4_port, QN => n_4632);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => n291, Q => 
                           REGISTERS_5_3_port, QN => n_4633);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => n361, Q => 
                           REGISTERS_5_2_port, QN => n_4634);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => n288, Q => 
                           REGISTERS_5_1_port, QN => n_4635);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => n368, Q => 
                           REGISTERS_5_0_port, QN => n_4636);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => n371, Q => 
                           REGISTERS_6_31_port, QN => n_4637);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => n374, Q => 
                           REGISTERS_6_30_port, QN => n_4638);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => n377, Q => 
                           REGISTERS_6_29_port, QN => n_4639);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => n380, Q => 
                           REGISTERS_6_28_port, QN => n_4640);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => n383, Q => 
                           REGISTERS_6_27_port, QN => n_4641);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => n365, Q => 
                           REGISTERS_6_26_port, QN => n_4642);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => n352, Q => 
                           REGISTERS_6_25_port, QN => n_4643);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => n355, Q => 
                           REGISTERS_6_24_port, QN => n_4644);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => n343, Q => 
                           REGISTERS_6_23_port, QN => n_4645);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => n346, Q => 
                           REGISTERS_6_22_port, QN => n_4646);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => n349, Q => 
                           REGISTERS_6_21_port, QN => n_4647);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => n331, Q => 
                           REGISTERS_6_20_port, QN => n_4648);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => n334, Q => 
                           REGISTERS_6_19_port, QN => n_4649);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => n337, Q => 
                           REGISTERS_6_18_port, QN => n_4650);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => n358, Q => 
                           REGISTERS_6_17_port, QN => n_4651);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => n340, Q => 
                           REGISTERS_6_16_port, QN => n_4652);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => n325, Q => 
                           REGISTERS_6_15_port, QN => n_4653);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => n328, Q => 
                           REGISTERS_6_14_port, QN => n_4654);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => n322, Q => 
                           REGISTERS_6_13_port, QN => n_4655);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => n319, Q => 
                           REGISTERS_6_12_port, QN => n_4656);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => n315, Q => 
                           REGISTERS_6_11_port, QN => n_4657);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => n312, Q => 
                           REGISTERS_6_10_port, QN => n_4658);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => n309, Q => 
                           REGISTERS_6_9_port, QN => n_4659);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => n306, Q => 
                           REGISTERS_6_8_port, QN => n_4660);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => n303, Q => 
                           REGISTERS_6_7_port, QN => n_4661);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => n300, Q => 
                           REGISTERS_6_6_port, QN => n_4662);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => n297, Q => 
                           REGISTERS_6_5_port, QN => n_4663);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => n294, Q => 
                           REGISTERS_6_4_port, QN => n_4664);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => n291, Q => 
                           REGISTERS_6_3_port, QN => n_4665);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => n362, Q => 
                           REGISTERS_6_2_port, QN => n_4666);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => n288, Q => 
                           REGISTERS_6_1_port, QN => n_4667);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => n368, Q => 
                           REGISTERS_6_0_port, QN => n_4668);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => n371, Q => 
                           REGISTERS_7_31_port, QN => n_4669);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => n374, Q => 
                           REGISTERS_7_30_port, QN => n_4670);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => n377, Q => 
                           REGISTERS_7_29_port, QN => n_4671);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => n380, Q => 
                           REGISTERS_7_28_port, QN => n_4672);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => n383, Q => 
                           REGISTERS_7_27_port, QN => n_4673);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => n365, Q => 
                           REGISTERS_7_26_port, QN => n_4674);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => n352, Q => 
                           REGISTERS_7_25_port, QN => n_4675);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => n355, Q => 
                           REGISTERS_7_24_port, QN => n_4676);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => n343, Q => 
                           REGISTERS_7_23_port, QN => n_4677);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => n346, Q => 
                           REGISTERS_7_22_port, QN => n_4678);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => n349, Q => 
                           REGISTERS_7_21_port, QN => n_4679);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => n331, Q => 
                           REGISTERS_7_20_port, QN => n_4680);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => n334, Q => 
                           REGISTERS_7_19_port, QN => n_4681);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => n337, Q => 
                           REGISTERS_7_18_port, QN => n_4682);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => n359, Q => 
                           REGISTERS_7_17_port, QN => n_4683);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => n340, Q => 
                           REGISTERS_7_16_port, QN => n_4684);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => n325, Q => 
                           REGISTERS_7_15_port, QN => n_4685);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => n328, Q => 
                           REGISTERS_7_14_port, QN => n_4686);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => n322, Q => 
                           REGISTERS_7_13_port, QN => n_4687);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => n319, Q => 
                           REGISTERS_7_12_port, QN => n_4688);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => n316, Q => 
                           REGISTERS_7_11_port, QN => n_4689);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => n312, Q => 
                           REGISTERS_7_10_port, QN => n_4690);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => n309, Q => 
                           REGISTERS_7_9_port, QN => n_4691);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => n306, Q => 
                           REGISTERS_7_8_port, QN => n_4692);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => n303, Q => 
                           REGISTERS_7_7_port, QN => n_4693);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => n300, Q => 
                           REGISTERS_7_6_port, QN => n_4694);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => n297, Q => 
                           REGISTERS_7_5_port, QN => n_4695);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => n294, Q => 
                           REGISTERS_7_4_port, QN => n_4696);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => n291, Q => 
                           REGISTERS_7_3_port, QN => n_4697);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => n362, Q => 
                           REGISTERS_7_2_port, QN => n_4698);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => n288, Q => 
                           REGISTERS_7_1_port, QN => n_4699);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => n368, Q => 
                           REGISTERS_7_0_port, QN => n_4700);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => n371, Q => 
                           REGISTERS_8_31_port, QN => n_4701);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => n374, Q => 
                           REGISTERS_8_30_port, QN => n_4702);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => n377, Q => 
                           REGISTERS_8_29_port, QN => n_4703);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => n380, Q => 
                           REGISTERS_8_28_port, QN => n_4704);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => n383, Q => 
                           REGISTERS_8_27_port, QN => n_4705);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => n365, Q => 
                           REGISTERS_8_26_port, QN => n_4706);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => n352, Q => 
                           REGISTERS_8_25_port, QN => n_4707);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => n356, Q => 
                           REGISTERS_8_24_port, QN => n_4708);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => n343, Q => 
                           REGISTERS_8_23_port, QN => n_4709);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => n346, Q => 
                           REGISTERS_8_22_port, QN => n_4710);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => n349, Q => 
                           REGISTERS_8_21_port, QN => n_4711);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => n331, Q => 
                           REGISTERS_8_20_port, QN => n_4712);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => n334, Q => 
                           REGISTERS_8_19_port, QN => n_4713);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => n337, Q => 
                           REGISTERS_8_18_port, QN => n_4714);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => n359, Q => 
                           REGISTERS_8_17_port, QN => n_4715);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => n340, Q => 
                           REGISTERS_8_16_port, QN => n_4716);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => n325, Q => 
                           REGISTERS_8_15_port, QN => n_4717);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => n328, Q => 
                           REGISTERS_8_14_port, QN => n_4718);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => n322, Q => 
                           REGISTERS_8_13_port, QN => n_4719);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => n319, Q => 
                           REGISTERS_8_12_port, QN => n_4720);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => n316, Q => 
                           REGISTERS_8_11_port, QN => n_4721);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => n313, Q => 
                           REGISTERS_8_10_port, QN => n_4722);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => n309, Q => 
                           REGISTERS_8_9_port, QN => n_4723);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => n306, Q => 
                           REGISTERS_8_8_port, QN => n_4724);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => n303, Q => 
                           REGISTERS_8_7_port, QN => n_4725);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => n300, Q => 
                           REGISTERS_8_6_port, QN => n_4726);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => n297, Q => 
                           REGISTERS_8_5_port, QN => n_4727);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => n294, Q => 
                           REGISTERS_8_4_port, QN => n_4728);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => n291, Q => 
                           REGISTERS_8_3_port, QN => n_4729);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => n362, Q => 
                           REGISTERS_8_2_port, QN => n_4730);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => n288, Q => 
                           REGISTERS_8_1_port, QN => n_4731);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => n368, Q => 
                           REGISTERS_8_0_port, QN => n_4732);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => n371, Q => 
                           REGISTERS_9_31_port, QN => n_4733);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => n374, Q => 
                           REGISTERS_9_30_port, QN => n_4734);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => n377, Q => 
                           REGISTERS_9_29_port, QN => n_4735);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => n380, Q => 
                           REGISTERS_9_28_port, QN => n_4736);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => n383, Q => 
                           REGISTERS_9_27_port, QN => n_4737);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => n365, Q => 
                           REGISTERS_9_26_port, QN => n_4738);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => n353, Q => 
                           REGISTERS_9_25_port, QN => n_4739);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => n356, Q => 
                           REGISTERS_9_24_port, QN => n_4740);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => n343, Q => 
                           REGISTERS_9_23_port, QN => n_4741);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => n346, Q => 
                           REGISTERS_9_22_port, QN => n_4742);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => n350, Q => 
                           REGISTERS_9_21_port, QN => n_4743);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => n331, Q => 
                           REGISTERS_9_20_port, QN => n_4744);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => n334, Q => 
                           REGISTERS_9_19_port, QN => n_4745);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => n337, Q => 
                           REGISTERS_9_18_port, QN => n_4746);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => n359, Q => 
                           REGISTERS_9_17_port, QN => n_4747);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => n340, Q => 
                           REGISTERS_9_16_port, QN => n_4748);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => n325, Q => 
                           REGISTERS_9_15_port, QN => n_4749);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => n328, Q => 
                           REGISTERS_9_14_port, QN => n_4750);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => n322, Q => 
                           REGISTERS_9_13_port, QN => n_4751);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => n319, Q => 
                           REGISTERS_9_12_port, QN => n_4752);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => n316, Q => 
                           REGISTERS_9_11_port, QN => n_4753);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => n313, Q => 
                           REGISTERS_9_10_port, QN => n_4754);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => n310, Q => 
                           REGISTERS_9_9_port, QN => n_4755);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => n306, Q => 
                           REGISTERS_9_8_port, QN => n_4756);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => n303, Q => 
                           REGISTERS_9_7_port, QN => n_4757);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => n300, Q => 
                           REGISTERS_9_6_port, QN => n_4758);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => n297, Q => 
                           REGISTERS_9_5_port, QN => n_4759);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => n294, Q => 
                           REGISTERS_9_4_port, QN => n_4760);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => n291, Q => 
                           REGISTERS_9_3_port, QN => n_4761);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => n362, Q => 
                           REGISTERS_9_2_port, QN => n_4762);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => n288, Q => 
                           REGISTERS_9_1_port, QN => n_4763);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => n368, Q => 
                           REGISTERS_9_0_port, QN => n_4764);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => n371, Q => 
                           REGISTERS_10_31_port, QN => n_4765);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => n374, Q => 
                           REGISTERS_10_30_port, QN => n_4766);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => n377, Q => 
                           REGISTERS_10_29_port, QN => n_4767);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => n380, Q => 
                           REGISTERS_10_28_port, QN => n_4768);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => n383, Q => 
                           REGISTERS_10_27_port, QN => n_4769);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => n365, Q => 
                           REGISTERS_10_26_port, QN => n_4770);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => n353, Q => 
                           REGISTERS_10_25_port, QN => n_4771);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => n356, Q => 
                           REGISTERS_10_24_port, QN => n_4772);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => n343, Q => 
                           REGISTERS_10_23_port, QN => n_4773);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => n347, Q => 
                           REGISTERS_10_22_port, QN => n_4774);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => n350, Q => 
                           REGISTERS_10_21_port, QN => n_4775);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => n331, Q => 
                           REGISTERS_10_20_port, QN => n_4776);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => n334, Q => 
                           REGISTERS_10_19_port, QN => n_4777);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => n337, Q => 
                           REGISTERS_10_18_port, QN => n_4778);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => n359, Q => 
                           REGISTERS_10_17_port, QN => n_4779);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => n340, Q => 
                           REGISTERS_10_16_port, QN => n_4780);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => n325, Q => 
                           REGISTERS_10_15_port, QN => n_4781);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => n328, Q => 
                           REGISTERS_10_14_port, QN => n_4782);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => n322, Q => 
                           REGISTERS_10_13_port, QN => n_4783);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => n319, Q => 
                           REGISTERS_10_12_port, QN => n_4784);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => n316, Q => 
                           REGISTERS_10_11_port, QN => n_4785);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => n313, Q => 
                           REGISTERS_10_10_port, QN => n_4786);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => n310, Q => 
                           REGISTERS_10_9_port, QN => n_4787);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => n307, Q => 
                           REGISTERS_10_8_port, QN => n_4788);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => n303, Q => 
                           REGISTERS_10_7_port, QN => n_4789);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => n300, Q => 
                           REGISTERS_10_6_port, QN => n_4790);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => n297, Q => 
                           REGISTERS_10_5_port, QN => n_4791);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => n294, Q => 
                           REGISTERS_10_4_port, QN => n_4792);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => n291, Q => 
                           REGISTERS_10_3_port, QN => n_4793);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => n362, Q => 
                           REGISTERS_10_2_port, QN => n_4794);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => n288, Q => 
                           REGISTERS_10_1_port, QN => n_4795);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => n368, Q => 
                           REGISTERS_10_0_port, QN => n_4796);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => n371, Q => 
                           REGISTERS_11_31_port, QN => n_4797);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => n374, Q => 
                           REGISTERS_11_30_port, QN => n_4798);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => n377, Q => 
                           REGISTERS_11_29_port, QN => n_4799);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => n380, Q => 
                           REGISTERS_11_28_port, QN => n_4800);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => n384, Q => 
                           REGISTERS_11_27_port, QN => n_4801);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => n365, Q => 
                           REGISTERS_11_26_port, QN => n_4802);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => n353, Q => 
                           REGISTERS_11_25_port, QN => n_4803);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => n356, Q => 
                           REGISTERS_11_24_port, QN => n_4804);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => n344, Q => 
                           REGISTERS_11_23_port, QN => n_4805);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => n347, Q => 
                           REGISTERS_11_22_port, QN => n_4806);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => n350, Q => 
                           REGISTERS_11_21_port, QN => n_4807);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => n331, Q => 
                           REGISTERS_11_20_port, QN => n_4808);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => n334, Q => 
                           REGISTERS_11_19_port, QN => n_4809);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => n337, Q => 
                           REGISTERS_11_18_port, QN => n_4810);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => n359, Q => 
                           REGISTERS_11_17_port, QN => n_4811);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => n341, Q => 
                           REGISTERS_11_16_port, QN => n_4812);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => n325, Q => 
                           REGISTERS_11_15_port, QN => n_4813);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => n328, Q => 
                           REGISTERS_11_14_port, QN => n_4814);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => n322, Q => 
                           REGISTERS_11_13_port, QN => n_4815);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => n319, Q => 
                           REGISTERS_11_12_port, QN => n_4816);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => n316, Q => 
                           REGISTERS_11_11_port, QN => n_4817);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => n313, Q => 
                           REGISTERS_11_10_port, QN => n_4818);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => n310, Q => 
                           REGISTERS_11_9_port, QN => n_4819);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => n307, Q => 
                           REGISTERS_11_8_port, QN => n_4820);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => n304, Q => 
                           REGISTERS_11_7_port, QN => n_4821);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => n300, Q => 
                           REGISTERS_11_6_port, QN => n_4822);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => n297, Q => 
                           REGISTERS_11_5_port, QN => n_4823);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => n294, Q => 
                           REGISTERS_11_4_port, QN => n_4824);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => n291, Q => 
                           REGISTERS_11_3_port, QN => n_4825);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => n362, Q => 
                           REGISTERS_11_2_port, QN => n_4826);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => n288, Q => 
                           REGISTERS_11_1_port, QN => n_4827);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => n368, Q => 
                           REGISTERS_11_0_port, QN => n_4828);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => n371, Q => 
                           REGISTERS_12_31_port, QN => n_4829);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => n374, Q => 
                           REGISTERS_12_30_port, QN => n_4830);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => n377, Q => 
                           REGISTERS_12_29_port, QN => n_4831);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => n381, Q => 
                           REGISTERS_12_28_port, QN => n_4832);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => n384, Q => 
                           REGISTERS_12_27_port, QN => n_4833);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => n365, Q => 
                           REGISTERS_12_26_port, QN => n_4834);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => n353, Q => 
                           REGISTERS_12_25_port, QN => n_4835);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => n356, Q => 
                           REGISTERS_12_24_port, QN => n_4836);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => n344, Q => 
                           REGISTERS_12_23_port, QN => n_4837);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => n347, Q => 
                           REGISTERS_12_22_port, QN => n_4838);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => n350, Q => 
                           REGISTERS_12_21_port, QN => n_4839);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => n331, Q => 
                           REGISTERS_12_20_port, QN => n_4840);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => n334, Q => 
                           REGISTERS_12_19_port, QN => n_4841);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => n338, Q => 
                           REGISTERS_12_18_port, QN => n_4842);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => n359, Q => 
                           REGISTERS_12_17_port, QN => n_4843);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => n341, Q => 
                           REGISTERS_12_16_port, QN => n_4844);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => n325, Q => 
                           REGISTERS_12_15_port, QN => n_4845);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => n328, Q => 
                           REGISTERS_12_14_port, QN => n_4846);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => n322, Q => 
                           REGISTERS_12_13_port, QN => n_4847);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => n319, Q => 
                           REGISTERS_12_12_port, QN => n_4848);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => n316, Q => 
                           REGISTERS_12_11_port, QN => n_4849);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => n313, Q => 
                           REGISTERS_12_10_port, QN => n_4850);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => n310, Q => 
                           REGISTERS_12_9_port, QN => n_4851);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => n307, Q => 
                           REGISTERS_12_8_port, QN => n_4852);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => n304, Q => 
                           REGISTERS_12_7_port, QN => n_4853);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => n301, Q => 
                           REGISTERS_12_6_port, QN => n_4854);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => n297, Q => 
                           REGISTERS_12_5_port, QN => n_4855);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => n294, Q => 
                           REGISTERS_12_4_port, QN => n_4856);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => n291, Q => 
                           REGISTERS_12_3_port, QN => n_4857);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => n362, Q => 
                           REGISTERS_12_2_port, QN => n_4858);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => n288, Q => 
                           REGISTERS_12_1_port, QN => n_4859);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => n368, Q => 
                           REGISTERS_12_0_port, QN => n_4860);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => n371, Q => 
                           REGISTERS_13_31_port, QN => n_4861);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => n374, Q => 
                           REGISTERS_13_30_port, QN => n_4862);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => n378, Q => 
                           REGISTERS_13_29_port, QN => n_4863);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => n381, Q => 
                           REGISTERS_13_28_port, QN => n_4864);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => n384, Q => 
                           REGISTERS_13_27_port, QN => n_4865);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => n365, Q => 
                           REGISTERS_13_26_port, QN => n_4866);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => n353, Q => 
                           REGISTERS_13_25_port, QN => n_4867);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => n356, Q => 
                           REGISTERS_13_24_port, QN => n_4868);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => n344, Q => 
                           REGISTERS_13_23_port, QN => n_4869);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => n347, Q => 
                           REGISTERS_13_22_port, QN => n_4870);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => n350, Q => 
                           REGISTERS_13_21_port, QN => n_4871);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => n331, Q => 
                           REGISTERS_13_20_port, QN => n_4872);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => n335, Q => 
                           REGISTERS_13_19_port, QN => n_4873);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => n338, Q => 
                           REGISTERS_13_18_port, QN => n_4874);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => n359, Q => 
                           REGISTERS_13_17_port, QN => n_4875);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => n341, Q => 
                           REGISTERS_13_16_port, QN => n_4876);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => n325, Q => 
                           REGISTERS_13_15_port, QN => n_4877);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => n328, Q => 
                           REGISTERS_13_14_port, QN => n_4878);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => n322, Q => 
                           REGISTERS_13_13_port, QN => n_4879);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => n319, Q => 
                           REGISTERS_13_12_port, QN => n_4880);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => n316, Q => 
                           REGISTERS_13_11_port, QN => n_4881);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => n313, Q => 
                           REGISTERS_13_10_port, QN => n_4882);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => n310, Q => 
                           REGISTERS_13_9_port, QN => n_4883);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => n307, Q => 
                           REGISTERS_13_8_port, QN => n_4884);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => n304, Q => 
                           REGISTERS_13_7_port, QN => n_4885);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => n301, Q => 
                           REGISTERS_13_6_port, QN => n_4886);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => n298, Q => 
                           REGISTERS_13_5_port, QN => n_4887);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => n294, Q => 
                           REGISTERS_13_4_port, QN => n_4888);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => n291, Q => 
                           REGISTERS_13_3_port, QN => n_4889);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => n362, Q => 
                           REGISTERS_13_2_port, QN => n_4890);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => n288, Q => 
                           REGISTERS_13_1_port, QN => n_4891);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => n368, Q => 
                           REGISTERS_13_0_port, QN => n_4892);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => n371, Q => 
                           REGISTERS_14_31_port, QN => n_4893);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => n375, Q => 
                           REGISTERS_14_30_port, QN => n_4894);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => n378, Q => 
                           REGISTERS_14_29_port, QN => n_4895);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => n381, Q => 
                           REGISTERS_14_28_port, QN => n_4896);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => n384, Q => 
                           REGISTERS_14_27_port, QN => n_4897);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => n365, Q => 
                           REGISTERS_14_26_port, QN => n_4898);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => n353, Q => 
                           REGISTERS_14_25_port, QN => n_4899);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => n356, Q => 
                           REGISTERS_14_24_port, QN => n_4900);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => n344, Q => 
                           REGISTERS_14_23_port, QN => n_4901);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => n347, Q => 
                           REGISTERS_14_22_port, QN => n_4902);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => n350, Q => 
                           REGISTERS_14_21_port, QN => n_4903);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => n332, Q => 
                           REGISTERS_14_20_port, QN => n_4904);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => n335, Q => 
                           REGISTERS_14_19_port, QN => n_4905);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => n338, Q => 
                           REGISTERS_14_18_port, QN => n_4906);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => n359, Q => 
                           REGISTERS_14_17_port, QN => n_4907);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => n341, Q => 
                           REGISTERS_14_16_port, QN => n_4908);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => n325, Q => 
                           REGISTERS_14_15_port, QN => n_4909);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => n329, Q => 
                           REGISTERS_14_14_port, QN => n_4910);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => n322, Q => 
                           REGISTERS_14_13_port, QN => n_4911);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => n319, Q => 
                           REGISTERS_14_12_port, QN => n_4912);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => n316, Q => 
                           REGISTERS_14_11_port, QN => n_4913);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => n313, Q => 
                           REGISTERS_14_10_port, QN => n_4914);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => n310, Q => 
                           REGISTERS_14_9_port, QN => n_4915);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => n307, Q => 
                           REGISTERS_14_8_port, QN => n_4916);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => n304, Q => 
                           REGISTERS_14_7_port, QN => n_4917);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => n301, Q => 
                           REGISTERS_14_6_port, QN => n_4918);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => n298, Q => 
                           REGISTERS_14_5_port, QN => n_4919);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => n295, Q => 
                           REGISTERS_14_4_port, QN => n_4920);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => n291, Q => 
                           REGISTERS_14_3_port, QN => n_4921);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => n362, Q => 
                           REGISTERS_14_2_port, QN => n_4922);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => n288, Q => 
                           REGISTERS_14_1_port, QN => n_4923);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => n368, Q => 
                           REGISTERS_14_0_port, QN => n_4924);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => n372, Q => 
                           REGISTERS_15_31_port, QN => n_4925);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => n375, Q => 
                           REGISTERS_15_30_port, QN => n_4926);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => n378, Q => 
                           REGISTERS_15_29_port, QN => n_4927);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => n381, Q => 
                           REGISTERS_15_28_port, QN => n_4928);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => n384, Q => 
                           REGISTERS_15_27_port, QN => n_4929);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => n365, Q => 
                           REGISTERS_15_26_port, QN => n_4930);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => n353, Q => 
                           REGISTERS_15_25_port, QN => n_4931);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => n356, Q => 
                           REGISTERS_15_24_port, QN => n_4932);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => n344, Q => 
                           REGISTERS_15_23_port, QN => n_4933);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => n347, Q => 
                           REGISTERS_15_22_port, QN => n_4934);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => n350, Q => 
                           REGISTERS_15_21_port, QN => n_4935);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => n332, Q => 
                           REGISTERS_15_20_port, QN => n_4936);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => n335, Q => 
                           REGISTERS_15_19_port, QN => n_4937);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => n338, Q => 
                           REGISTERS_15_18_port, QN => n_4938);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => n359, Q => 
                           REGISTERS_15_17_port, QN => n_4939);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => n341, Q => 
                           REGISTERS_15_16_port, QN => n_4940);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => n326, Q => 
                           REGISTERS_15_15_port, QN => n_4941);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => n329, Q => 
                           REGISTERS_15_14_port, QN => n_4942);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => n322, Q => 
                           REGISTERS_15_13_port, QN => n_4943);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => n319, Q => 
                           REGISTERS_15_12_port, QN => n_4944);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => n316, Q => 
                           REGISTERS_15_11_port, QN => n_4945);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => n313, Q => 
                           REGISTERS_15_10_port, QN => n_4946);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => n310, Q => 
                           REGISTERS_15_9_port, QN => n_4947);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => n307, Q => 
                           REGISTERS_15_8_port, QN => n_4948);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => n304, Q => 
                           REGISTERS_15_7_port, QN => n_4949);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => n301, Q => 
                           REGISTERS_15_6_port, QN => n_4950);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => n298, Q => 
                           REGISTERS_15_5_port, QN => n_4951);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => n295, Q => 
                           REGISTERS_15_4_port, QN => n_4952);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => n292, Q => 
                           REGISTERS_15_3_port, QN => n_4953);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => n362, Q => 
                           REGISTERS_15_2_port, QN => n_4954);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => n288, Q => 
                           REGISTERS_15_1_port, QN => n_4955);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => n368, Q => 
                           REGISTERS_15_0_port, QN => n_4956);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => n372, Q => 
                           REGISTERS_16_31_port, QN => n_4957);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => n375, Q => 
                           REGISTERS_16_30_port, QN => n_4958);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => n378, Q => 
                           REGISTERS_16_29_port, QN => n_4959);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => n381, Q => 
                           REGISTERS_16_28_port, QN => n_4960);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => n384, Q => 
                           REGISTERS_16_27_port, QN => n_4961);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => n365, Q => 
                           REGISTERS_16_26_port, QN => n_4962);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => n353, Q => 
                           REGISTERS_16_25_port, QN => n_4963);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => n356, Q => 
                           REGISTERS_16_24_port, QN => n_4964);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => n344, Q => 
                           REGISTERS_16_23_port, QN => n_4965);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => n347, Q => 
                           REGISTERS_16_22_port, QN => n_4966);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => n350, Q => 
                           REGISTERS_16_21_port, QN => n_4967);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => n332, Q => 
                           REGISTERS_16_20_port, QN => n_4968);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => n335, Q => 
                           REGISTERS_16_19_port, QN => n_4969);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => n338, Q => 
                           REGISTERS_16_18_port, QN => n_4970);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => n359, Q => 
                           REGISTERS_16_17_port, QN => n_4971);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => n341, Q => 
                           REGISTERS_16_16_port, QN => n_4972);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => n326, Q => 
                           REGISTERS_16_15_port, QN => n_4973);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => n329, Q => 
                           REGISTERS_16_14_port, QN => n_4974);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => n323, Q => 
                           REGISTERS_16_13_port, QN => n_4975);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => n319, Q => 
                           REGISTERS_16_12_port, QN => n_4976);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => n316, Q => 
                           REGISTERS_16_11_port, QN => n_4977);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => n313, Q => 
                           REGISTERS_16_10_port, QN => n_4978);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => n310, Q => 
                           REGISTERS_16_9_port, QN => n_4979);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => n307, Q => 
                           REGISTERS_16_8_port, QN => n_4980);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => n304, Q => 
                           REGISTERS_16_7_port, QN => n_4981);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => n301, Q => 
                           REGISTERS_16_6_port, QN => n_4982);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => n298, Q => 
                           REGISTERS_16_5_port, QN => n_4983);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => n295, Q => 
                           REGISTERS_16_4_port, QN => n_4984);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => n292, Q => 
                           REGISTERS_16_3_port, QN => n_4985);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => n362, Q => 
                           REGISTERS_16_2_port, QN => n_4986);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => n289, Q => 
                           REGISTERS_16_1_port, QN => n_4987);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => n369, Q => 
                           REGISTERS_16_0_port, QN => n_4988);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => n372, Q => 
                           REGISTERS_17_31_port, QN => n_4989);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => n375, Q => 
                           REGISTERS_17_30_port, QN => n_4990);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => n378, Q => 
                           REGISTERS_17_29_port, QN => n_4991);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => n381, Q => 
                           REGISTERS_17_28_port, QN => n_4992);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => n384, Q => 
                           REGISTERS_17_27_port, QN => n_4993);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => n366, Q => 
                           REGISTERS_17_26_port, QN => n_4994);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => n353, Q => 
                           REGISTERS_17_25_port, QN => n_4995);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => n356, Q => 
                           REGISTERS_17_24_port, QN => n_4996);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => n344, Q => 
                           REGISTERS_17_23_port, QN => n_4997);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => n347, Q => 
                           REGISTERS_17_22_port, QN => n_4998);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => n350, Q => 
                           REGISTERS_17_21_port, QN => n_4999);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => n332, Q => 
                           REGISTERS_17_20_port, QN => n_5000);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => n335, Q => 
                           REGISTERS_17_19_port, QN => n_5001);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => n338, Q => 
                           REGISTERS_17_18_port, QN => n_5002);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => n359, Q => 
                           REGISTERS_17_17_port, QN => n_5003);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => n341, Q => 
                           REGISTERS_17_16_port, QN => n_5004);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => n326, Q => 
                           REGISTERS_17_15_port, QN => n_5005);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => n329, Q => 
                           REGISTERS_17_14_port, QN => n_5006);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => n323, Q => 
                           REGISTERS_17_13_port, QN => n_5007);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => n320, Q => 
                           REGISTERS_17_12_port, QN => n_5008);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => n316, Q => 
                           REGISTERS_17_11_port, QN => n_5009);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => n313, Q => 
                           REGISTERS_17_10_port, QN => n_5010);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => n310, Q => 
                           REGISTERS_17_9_port, QN => n_5011);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => n307, Q => 
                           REGISTERS_17_8_port, QN => n_5012);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => n304, Q => 
                           REGISTERS_17_7_port, QN => n_5013);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => n301, Q => 
                           REGISTERS_17_6_port, QN => n_5014);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => n298, Q => 
                           REGISTERS_17_5_port, QN => n_5015);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => n295, Q => 
                           REGISTERS_17_4_port, QN => n_5016);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => n292, Q => 
                           REGISTERS_17_3_port, QN => n_5017);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => n363, Q => 
                           REGISTERS_17_2_port, QN => n_5018);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => n289, Q => 
                           REGISTERS_17_1_port, QN => n_5019);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => n369, Q => 
                           REGISTERS_17_0_port, QN => n_5020);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => n372, Q => 
                           REGISTERS_18_31_port, QN => n_5021);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => n375, Q => 
                           REGISTERS_18_30_port, QN => n_5022);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => n378, Q => 
                           REGISTERS_18_29_port, QN => n_5023);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => n381, Q => 
                           REGISTERS_18_28_port, QN => n_5024);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => n384, Q => 
                           REGISTERS_18_27_port, QN => n_5025);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => n366, Q => 
                           REGISTERS_18_26_port, QN => n_5026);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => n353, Q => 
                           REGISTERS_18_25_port, QN => n_5027);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => n356, Q => 
                           REGISTERS_18_24_port, QN => n_5028);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => n344, Q => 
                           REGISTERS_18_23_port, QN => n_5029);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => n347, Q => 
                           REGISTERS_18_22_port, QN => n_5030);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => n350, Q => 
                           REGISTERS_18_21_port, QN => n_5031);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => n332, Q => 
                           REGISTERS_18_20_port, QN => n_5032);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => n335, Q => 
                           REGISTERS_18_19_port, QN => n_5033);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => n338, Q => 
                           REGISTERS_18_18_port, QN => n_5034);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => n360, Q => 
                           REGISTERS_18_17_port, QN => n_5035);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => n341, Q => 
                           REGISTERS_18_16_port, QN => n_5036);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => n326, Q => 
                           REGISTERS_18_15_port, QN => n_5037);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => n329, Q => 
                           REGISTERS_18_14_port, QN => n_5038);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => n323, Q => 
                           REGISTERS_18_13_port, QN => n_5039);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => n320, Q => 
                           REGISTERS_18_12_port, QN => n_5040);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => n317, Q => 
                           REGISTERS_18_11_port, QN => n_5041);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => n313, Q => 
                           REGISTERS_18_10_port, QN => n_5042);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => n310, Q => 
                           REGISTERS_18_9_port, QN => n_5043);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => n307, Q => 
                           REGISTERS_18_8_port, QN => n_5044);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => n304, Q => 
                           REGISTERS_18_7_port, QN => n_5045);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => n301, Q => 
                           REGISTERS_18_6_port, QN => n_5046);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => n298, Q => 
                           REGISTERS_18_5_port, QN => n_5047);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => n295, Q => 
                           REGISTERS_18_4_port, QN => n_5048);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => n292, Q => 
                           REGISTERS_18_3_port, QN => n_5049);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => n363, Q => 
                           REGISTERS_18_2_port, QN => n_5050);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => n289, Q => 
                           REGISTERS_18_1_port, QN => n_5051);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => n369, Q => 
                           REGISTERS_18_0_port, QN => n_5052);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => n372, Q => 
                           REGISTERS_19_31_port, QN => n_5053);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => n375, Q => 
                           REGISTERS_19_30_port, QN => n_5054);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => n378, Q => 
                           REGISTERS_19_29_port, QN => n_5055);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => n381, Q => 
                           REGISTERS_19_28_port, QN => n_5056);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => n384, Q => 
                           REGISTERS_19_27_port, QN => n_5057);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => n366, Q => 
                           REGISTERS_19_26_port, QN => n_5058);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => n353, Q => 
                           REGISTERS_19_25_port, QN => n_5059);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => n357, Q => 
                           REGISTERS_19_24_port, QN => n_5060);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => n344, Q => 
                           REGISTERS_19_23_port, QN => n_5061);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => n347, Q => 
                           REGISTERS_19_22_port, QN => n_5062);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => n350, Q => 
                           REGISTERS_19_21_port, QN => n_5063);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => n332, Q => 
                           REGISTERS_19_20_port, QN => n_5064);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => n335, Q => 
                           REGISTERS_19_19_port, QN => n_5065);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => n338, Q => 
                           REGISTERS_19_18_port, QN => n_5066);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => n360, Q => 
                           REGISTERS_19_17_port, QN => n_5067);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => n341, Q => 
                           REGISTERS_19_16_port, QN => n_5068);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => n326, Q => 
                           REGISTERS_19_15_port, QN => n_5069);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => n329, Q => 
                           REGISTERS_19_14_port, QN => n_5070);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => n323, Q => 
                           REGISTERS_19_13_port, QN => n_5071);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => n320, Q => 
                           REGISTERS_19_12_port, QN => n_5072);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => n317, Q => 
                           REGISTERS_19_11_port, QN => n_5073);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => n314, Q => 
                           REGISTERS_19_10_port, QN => n_5074);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => n310, Q => 
                           REGISTERS_19_9_port, QN => n_5075);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => n307, Q => 
                           REGISTERS_19_8_port, QN => n_5076);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => n304, Q => 
                           REGISTERS_19_7_port, QN => n_5077);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => n301, Q => 
                           REGISTERS_19_6_port, QN => n_5078);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => n298, Q => 
                           REGISTERS_19_5_port, QN => n_5079);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => n295, Q => 
                           REGISTERS_19_4_port, QN => n_5080);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => n292, Q => 
                           REGISTERS_19_3_port, QN => n_5081);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => n363, Q => 
                           REGISTERS_19_2_port, QN => n_5082);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => n289, Q => 
                           REGISTERS_19_1_port, QN => n_5083);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => n369, Q => 
                           REGISTERS_19_0_port, QN => n_5084);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => n372, Q => 
                           REGISTERS_20_31_port, QN => n_5085);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => n375, Q => 
                           REGISTERS_20_30_port, QN => n_5086);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => n378, Q => 
                           REGISTERS_20_29_port, QN => n_5087);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => n381, Q => 
                           REGISTERS_20_28_port, QN => n_5088);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => n384, Q => 
                           REGISTERS_20_27_port, QN => n_5089);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => n366, Q => 
                           REGISTERS_20_26_port, QN => n_5090);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => n354, Q => 
                           REGISTERS_20_25_port, QN => n_5091);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => n357, Q => 
                           REGISTERS_20_24_port, QN => n_5092);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => n344, Q => 
                           REGISTERS_20_23_port, QN => n_5093);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => n347, Q => 
                           REGISTERS_20_22_port, QN => n_5094);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => n351, Q => 
                           REGISTERS_20_21_port, QN => n_5095);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => n332, Q => 
                           REGISTERS_20_20_port, QN => n_5096);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => n335, Q => 
                           REGISTERS_20_19_port, QN => n_5097);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => n338, Q => 
                           REGISTERS_20_18_port, QN => n_5098);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => n360, Q => 
                           REGISTERS_20_17_port, QN => n_5099);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => n341, Q => 
                           REGISTERS_20_16_port, QN => n_5100);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => n326, Q => 
                           REGISTERS_20_15_port, QN => n_5101);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => n329, Q => 
                           REGISTERS_20_14_port, QN => n_5102);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => n323, Q => 
                           REGISTERS_20_13_port, QN => n_5103);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => n320, Q => 
                           REGISTERS_20_12_port, QN => n_5104);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => n317, Q => 
                           REGISTERS_20_11_port, QN => n_5105);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => n314, Q => 
                           REGISTERS_20_10_port, QN => n_5106);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => n311, Q => 
                           REGISTERS_20_9_port, QN => n_5107);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => n307, Q => 
                           REGISTERS_20_8_port, QN => n_5108);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => n304, Q => 
                           REGISTERS_20_7_port, QN => n_5109);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => n301, Q => 
                           REGISTERS_20_6_port, QN => n_5110);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => n298, Q => 
                           REGISTERS_20_5_port, QN => n_5111);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => n295, Q => 
                           REGISTERS_20_4_port, QN => n_5112);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => n292, Q => 
                           REGISTERS_20_3_port, QN => n_5113);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => n363, Q => 
                           REGISTERS_20_2_port, QN => n_5114);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => n289, Q => 
                           REGISTERS_20_1_port, QN => n_5115);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => n369, Q => 
                           REGISTERS_20_0_port, QN => n_5116);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => n372, Q => 
                           REGISTERS_21_31_port, QN => n_5117);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => n375, Q => 
                           REGISTERS_21_30_port, QN => n_5118);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => n378, Q => 
                           REGISTERS_21_29_port, QN => n_5119);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => n381, Q => 
                           REGISTERS_21_28_port, QN => n_5120);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => n384, Q => 
                           REGISTERS_21_27_port, QN => n_5121);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => n366, Q => 
                           REGISTERS_21_26_port, QN => n_5122);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => n354, Q => 
                           REGISTERS_21_25_port, QN => n_5123);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => n357, Q => 
                           REGISTERS_21_24_port, QN => n_5124);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => n344, Q => 
                           REGISTERS_21_23_port, QN => n_5125);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => n348, Q => 
                           REGISTERS_21_22_port, QN => n_5126);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => n351, Q => 
                           REGISTERS_21_21_port, QN => n_5127);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => n332, Q => 
                           REGISTERS_21_20_port, QN => n_5128);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => n335, Q => 
                           REGISTERS_21_19_port, QN => n_5129);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => n338, Q => 
                           REGISTERS_21_18_port, QN => n_5130);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => n360, Q => 
                           REGISTERS_21_17_port, QN => n_5131);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => n341, Q => 
                           REGISTERS_21_16_port, QN => n_5132);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => n326, Q => 
                           REGISTERS_21_15_port, QN => n_5133);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => n329, Q => 
                           REGISTERS_21_14_port, QN => n_5134);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => n323, Q => 
                           REGISTERS_21_13_port, QN => n_5135);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => n320, Q => 
                           REGISTERS_21_12_port, QN => n_5136);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => n317, Q => 
                           REGISTERS_21_11_port, QN => n_5137);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => n314, Q => 
                           REGISTERS_21_10_port, QN => n_5138);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => n311, Q => 
                           REGISTERS_21_9_port, QN => n_5139);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => n308, Q => 
                           REGISTERS_21_8_port, QN => n_5140);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => n304, Q => 
                           REGISTERS_21_7_port, QN => n_5141);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => n301, Q => 
                           REGISTERS_21_6_port, QN => n_5142);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => n298, Q => 
                           REGISTERS_21_5_port, QN => n_5143);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => n295, Q => 
                           REGISTERS_21_4_port, QN => n_5144);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => n292, Q => 
                           REGISTERS_21_3_port, QN => n_5145);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => n363, Q => 
                           REGISTERS_21_2_port, QN => n_5146);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => n289, Q => 
                           REGISTERS_21_1_port, QN => n_5147);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => n369, Q => 
                           REGISTERS_21_0_port, QN => n_5148);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => n372, Q => 
                           REGISTERS_22_31_port, QN => n_5149);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => n375, Q => 
                           REGISTERS_22_30_port, QN => n_5150);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => n378, Q => 
                           REGISTERS_22_29_port, QN => n_5151);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => n381, Q => 
                           REGISTERS_22_28_port, QN => n_5152);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => n385_port, Q 
                           => REGISTERS_22_27_port, QN => n_5153);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => n366, Q => 
                           REGISTERS_22_26_port, QN => n_5154);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => n354, Q => 
                           REGISTERS_22_25_port, QN => n_5155);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => n357, Q => 
                           REGISTERS_22_24_port, QN => n_5156);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => n345, Q => 
                           REGISTERS_22_23_port, QN => n_5157);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => n348, Q => 
                           REGISTERS_22_22_port, QN => n_5158);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => n351, Q => 
                           REGISTERS_22_21_port, QN => n_5159);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => n332, Q => 
                           REGISTERS_22_20_port, QN => n_5160);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => n335, Q => 
                           REGISTERS_22_19_port, QN => n_5161);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => n338, Q => 
                           REGISTERS_22_18_port, QN => n_5162);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => n360, Q => 
                           REGISTERS_22_17_port, QN => n_5163);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => n342, Q => 
                           REGISTERS_22_16_port, QN => n_5164);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => n326, Q => 
                           REGISTERS_22_15_port, QN => n_5165);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => n329, Q => 
                           REGISTERS_22_14_port, QN => n_5166);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => n323, Q => 
                           REGISTERS_22_13_port, QN => n_5167);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => n320, Q => 
                           REGISTERS_22_12_port, QN => n_5168);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => n317, Q => 
                           REGISTERS_22_11_port, QN => n_5169);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => n314, Q => 
                           REGISTERS_22_10_port, QN => n_5170);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => n311, Q => 
                           REGISTERS_22_9_port, QN => n_5171);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => n308, Q => 
                           REGISTERS_22_8_port, QN => n_5172);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => n305, Q => 
                           REGISTERS_22_7_port, QN => n_5173);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => n301, Q => 
                           REGISTERS_22_6_port, QN => n_5174);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => n298, Q => 
                           REGISTERS_22_5_port, QN => n_5175);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => n295, Q => 
                           REGISTERS_22_4_port, QN => n_5176);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => n292, Q => 
                           REGISTERS_22_3_port, QN => n_5177);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => n363, Q => 
                           REGISTERS_22_2_port, QN => n_5178);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => n289, Q => 
                           REGISTERS_22_1_port, QN => n_5179);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => n369, Q => 
                           REGISTERS_22_0_port, QN => n_5180);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => n372, Q => 
                           REGISTERS_23_31_port, QN => n_5181);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => n375, Q => 
                           REGISTERS_23_30_port, QN => n_5182);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => n378, Q => 
                           REGISTERS_23_29_port, QN => n_5183);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => n382, Q => 
                           REGISTERS_23_28_port, QN => n_5184);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => n385_port, Q 
                           => REGISTERS_23_27_port, QN => n_5185);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => n366, Q => 
                           REGISTERS_23_26_port, QN => n_5186);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => n354, Q => 
                           REGISTERS_23_25_port, QN => n_5187);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => n357, Q => 
                           REGISTERS_23_24_port, QN => n_5188);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => n345, Q => 
                           REGISTERS_23_23_port, QN => n_5189);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => n348, Q => 
                           REGISTERS_23_22_port, QN => n_5190);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => n351, Q => 
                           REGISTERS_23_21_port, QN => n_5191);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => n332, Q => 
                           REGISTERS_23_20_port, QN => n_5192);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => n335, Q => 
                           REGISTERS_23_19_port, QN => n_5193);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => n339, Q => 
                           REGISTERS_23_18_port, QN => n_5194);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => n360, Q => 
                           REGISTERS_23_17_port, QN => n_5195);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => n342, Q => 
                           REGISTERS_23_16_port, QN => n_5196);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => n326, Q => 
                           REGISTERS_23_15_port, QN => n_5197);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => n329, Q => 
                           REGISTERS_23_14_port, QN => n_5198);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => n323, Q => 
                           REGISTERS_23_13_port, QN => n_5199);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => n320, Q => 
                           REGISTERS_23_12_port, QN => n_5200);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => n317, Q => 
                           REGISTERS_23_11_port, QN => n_5201);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => n314, Q => 
                           REGISTERS_23_10_port, QN => n_5202);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => n311, Q => 
                           REGISTERS_23_9_port, QN => n_5203);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => n308, Q => 
                           REGISTERS_23_8_port, QN => n_5204);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => n305, Q => 
                           REGISTERS_23_7_port, QN => n_5205);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => n302, Q => 
                           REGISTERS_23_6_port, QN => n_5206);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => n298, Q => 
                           REGISTERS_23_5_port, QN => n_5207);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => n295, Q => 
                           REGISTERS_23_4_port, QN => n_5208);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => n292, Q => 
                           REGISTERS_23_3_port, QN => n_5209);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => n363, Q => 
                           REGISTERS_23_2_port, QN => n_5210);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => n289, Q => 
                           REGISTERS_23_1_port, QN => n_5211);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => n369, Q => 
                           REGISTERS_23_0_port, QN => n_5212);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => n372, Q => 
                           REGISTERS_24_31_port, QN => n_5213);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => n375, Q => 
                           REGISTERS_24_30_port, QN => n_5214);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => n379, Q => 
                           REGISTERS_24_29_port, QN => n_5215);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => n382, Q => 
                           REGISTERS_24_28_port, QN => n_5216);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => n385_port, Q 
                           => REGISTERS_24_27_port, QN => n_5217);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => n366, Q => 
                           REGISTERS_24_26_port, QN => n_5218);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => n354, Q => 
                           REGISTERS_24_25_port, QN => n_5219);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => n357, Q => 
                           REGISTERS_24_24_port, QN => n_5220);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => n345, Q => 
                           REGISTERS_24_23_port, QN => n_5221);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => n348, Q => 
                           REGISTERS_24_22_port, QN => n_5222);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => n351, Q => 
                           REGISTERS_24_21_port, QN => n_5223);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => n332, Q => 
                           REGISTERS_24_20_port, QN => n_5224);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => n336, Q => 
                           REGISTERS_24_19_port, QN => n_5225);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => n339, Q => 
                           REGISTERS_24_18_port, QN => n_5226);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => n360, Q => 
                           REGISTERS_24_17_port, QN => n_5227);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => n342, Q => 
                           REGISTERS_24_16_port, QN => n_5228);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => n326, Q => 
                           REGISTERS_24_15_port, QN => n_5229);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => n329, Q => 
                           REGISTERS_24_14_port, QN => n_5230);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => n323, Q => 
                           REGISTERS_24_13_port, QN => n_5231);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => n320, Q => 
                           REGISTERS_24_12_port, QN => n_5232);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => n317, Q => 
                           REGISTERS_24_11_port, QN => n_5233);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => n314, Q => 
                           REGISTERS_24_10_port, QN => n_5234);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => n311, Q => 
                           REGISTERS_24_9_port, QN => n_5235);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => n308, Q => 
                           REGISTERS_24_8_port, QN => n_5236);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => n305, Q => 
                           REGISTERS_24_7_port, QN => n_5237);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => n302, Q => 
                           REGISTERS_24_6_port, QN => n_5238);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => n299, Q => 
                           REGISTERS_24_5_port, QN => n_5239);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => n295, Q => 
                           REGISTERS_24_4_port, QN => n_5240);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => n292, Q => 
                           REGISTERS_24_3_port, QN => n_5241);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => n363, Q => 
                           REGISTERS_24_2_port, QN => n_5242);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => n289, Q => 
                           REGISTERS_24_1_port, QN => n_5243);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => n369, Q => 
                           REGISTERS_24_0_port, QN => n_5244);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => n372, Q => 
                           REGISTERS_25_31_port, QN => n_5245);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => n376, Q => 
                           REGISTERS_25_30_port, QN => n_5246);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => n379, Q => 
                           REGISTERS_25_29_port, QN => n_5247);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => n382, Q => 
                           REGISTERS_25_28_port, QN => n_5248);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => n385_port, Q 
                           => REGISTERS_25_27_port, QN => n_5249);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => n366, Q => 
                           REGISTERS_25_26_port, QN => n_5250);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => n354, Q => 
                           REGISTERS_25_25_port, QN => n_5251);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => n357, Q => 
                           REGISTERS_25_24_port, QN => n_5252);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => n345, Q => 
                           REGISTERS_25_23_port, QN => n_5253);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => n348, Q => 
                           REGISTERS_25_22_port, QN => n_5254);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => n351, Q => 
                           REGISTERS_25_21_port, QN => n_5255);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => n333, Q => 
                           REGISTERS_25_20_port, QN => n_5256);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => n336, Q => 
                           REGISTERS_25_19_port, QN => n_5257);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => n339, Q => 
                           REGISTERS_25_18_port, QN => n_5258);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => n360, Q => 
                           REGISTERS_25_17_port, QN => n_5259);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => n342, Q => 
                           REGISTERS_25_16_port, QN => n_5260);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => n326, Q => 
                           REGISTERS_25_15_port, QN => n_5261);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => n330, Q => 
                           REGISTERS_25_14_port, QN => n_5262);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => n323, Q => 
                           REGISTERS_25_13_port, QN => n_5263);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => n320, Q => 
                           REGISTERS_25_12_port, QN => n_5264);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => n317, Q => 
                           REGISTERS_25_11_port, QN => n_5265);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => n314, Q => 
                           REGISTERS_25_10_port, QN => n_5266);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => n311, Q => 
                           REGISTERS_25_9_port, QN => n_5267);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => n308, Q => 
                           REGISTERS_25_8_port, QN => n_5268);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => n305, Q => 
                           REGISTERS_25_7_port, QN => n_5269);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => n302, Q => 
                           REGISTERS_25_6_port, QN => n_5270);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => n299, Q => 
                           REGISTERS_25_5_port, QN => n_5271);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => n296, Q => 
                           REGISTERS_25_4_port, QN => n_5272);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => n292, Q => 
                           REGISTERS_25_3_port, QN => n_5273);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => n363, Q => 
                           REGISTERS_25_2_port, QN => n_5274);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => n289, Q => 
                           REGISTERS_25_1_port, QN => n_5275);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => n369, Q => 
                           REGISTERS_25_0_port, QN => n_5276);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => n373, Q => 
                           REGISTERS_26_31_port, QN => n_5277);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => n376, Q => 
                           REGISTERS_26_30_port, QN => n_5278);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => n379, Q => 
                           REGISTERS_26_29_port, QN => n_5279);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => n382, Q => 
                           REGISTERS_26_28_port, QN => n_5280);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => n385_port, Q 
                           => REGISTERS_26_27_port, QN => n_5281);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => n366, Q => 
                           REGISTERS_26_26_port, QN => n_5282);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => n354, Q => 
                           REGISTERS_26_25_port, QN => n_5283);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => n357, Q => 
                           REGISTERS_26_24_port, QN => n_5284);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => n345, Q => 
                           REGISTERS_26_23_port, QN => n_5285);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => n348, Q => 
                           REGISTERS_26_22_port, QN => n_5286);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => n351, Q => 
                           REGISTERS_26_21_port, QN => n_5287);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => n333, Q => 
                           REGISTERS_26_20_port, QN => n_5288);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => n336, Q => 
                           REGISTERS_26_19_port, QN => n_5289);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => n339, Q => 
                           REGISTERS_26_18_port, QN => n_5290);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => n360, Q => 
                           REGISTERS_26_17_port, QN => n_5291);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => n342, Q => 
                           REGISTERS_26_16_port, QN => n_5292);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => n327, Q => 
                           REGISTERS_26_15_port, QN => n_5293);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => n330, Q => 
                           REGISTERS_26_14_port, QN => n_5294);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => n323, Q => 
                           REGISTERS_26_13_port, QN => n_5295);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => n320, Q => 
                           REGISTERS_26_12_port, QN => n_5296);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => n317, Q => 
                           REGISTERS_26_11_port, QN => n_5297);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => n314, Q => 
                           REGISTERS_26_10_port, QN => n_5298);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => n311, Q => 
                           REGISTERS_26_9_port, QN => n_5299);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => n308, Q => 
                           REGISTERS_26_8_port, QN => n_5300);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => n305, Q => 
                           REGISTERS_26_7_port, QN => n_5301);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => n302, Q => 
                           REGISTERS_26_6_port, QN => n_5302);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => n299, Q => 
                           REGISTERS_26_5_port, QN => n_5303);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => n296, Q => 
                           REGISTERS_26_4_port, QN => n_5304);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => n293, Q => 
                           REGISTERS_26_3_port, QN => n_5305);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => n363, Q => 
                           REGISTERS_26_2_port, QN => n_5306);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => n289, Q => 
                           REGISTERS_26_1_port, QN => n_5307);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => n369, Q => 
                           REGISTERS_26_0_port, QN => n_5308);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => n373, Q => 
                           REGISTERS_27_31_port, QN => n_5309);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => n376, Q => 
                           REGISTERS_27_30_port, QN => n_5310);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => n379, Q => 
                           REGISTERS_27_29_port, QN => n_5311);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => n382, Q => 
                           REGISTERS_27_28_port, QN => n_5312);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => n385_port, Q 
                           => REGISTERS_27_27_port, QN => n_5313);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => n366, Q => 
                           REGISTERS_27_26_port, QN => n_5314);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => n354, Q => 
                           REGISTERS_27_25_port, QN => n_5315);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => n357, Q => 
                           REGISTERS_27_24_port, QN => n_5316);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => n345, Q => 
                           REGISTERS_27_23_port, QN => n_5317);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => n348, Q => 
                           REGISTERS_27_22_port, QN => n_5318);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => n351, Q => 
                           REGISTERS_27_21_port, QN => n_5319);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => n333, Q => 
                           REGISTERS_27_20_port, QN => n_5320);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => n336, Q => 
                           REGISTERS_27_19_port, QN => n_5321);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => n339, Q => 
                           REGISTERS_27_18_port, QN => n_5322);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => n360, Q => 
                           REGISTERS_27_17_port, QN => n_5323);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => n342, Q => 
                           REGISTERS_27_16_port, QN => n_5324);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => n327, Q => 
                           REGISTERS_27_15_port, QN => n_5325);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => n330, Q => 
                           REGISTERS_27_14_port, QN => n_5326);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => n324, Q => 
                           REGISTERS_27_13_port, QN => n_5327);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => n320, Q => 
                           REGISTERS_27_12_port, QN => n_5328);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => n317, Q => 
                           REGISTERS_27_11_port, QN => n_5329);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => n314, Q => 
                           REGISTERS_27_10_port, QN => n_5330);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => n311, Q => 
                           REGISTERS_27_9_port, QN => n_5331);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => n308, Q => 
                           REGISTERS_27_8_port, QN => n_5332);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => n305, Q => 
                           REGISTERS_27_7_port, QN => n_5333);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => n302, Q => 
                           REGISTERS_27_6_port, QN => n_5334);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => n299, Q => 
                           REGISTERS_27_5_port, QN => n_5335);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => n296, Q => 
                           REGISTERS_27_4_port, QN => n_5336);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => n293, Q => 
                           REGISTERS_27_3_port, QN => n_5337);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => n363, Q => 
                           REGISTERS_27_2_port, QN => n_5338);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => n290, Q => 
                           REGISTERS_27_1_port, QN => n_5339);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => n370, Q => 
                           REGISTERS_27_0_port, QN => n_5340);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => n373, Q => 
                           REGISTERS_28_31_port, QN => n_5341);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => n376, Q => 
                           REGISTERS_28_30_port, QN => n_5342);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => n379, Q => 
                           REGISTERS_28_29_port, QN => n_5343);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => n382, Q => 
                           REGISTERS_28_28_port, QN => n_5344);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => n385_port, Q 
                           => REGISTERS_28_27_port, QN => n_5345);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => n367, Q => 
                           REGISTERS_28_26_port, QN => n_5346);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => n354, Q => 
                           REGISTERS_28_25_port, QN => n_5347);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => n357, Q => 
                           REGISTERS_28_24_port, QN => n_5348);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => n345, Q => 
                           REGISTERS_28_23_port, QN => n_5349);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => n348, Q => 
                           REGISTERS_28_22_port, QN => n_5350);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => n351, Q => 
                           REGISTERS_28_21_port, QN => n_5351);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => n333, Q => 
                           REGISTERS_28_20_port, QN => n_5352);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => n336, Q => 
                           REGISTERS_28_19_port, QN => n_5353);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => n339, Q => 
                           REGISTERS_28_18_port, QN => n_5354);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => n360, Q => 
                           REGISTERS_28_17_port, QN => n_5355);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => n342, Q => 
                           REGISTERS_28_16_port, QN => n_5356);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => n327, Q => 
                           REGISTERS_28_15_port, QN => n_5357);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => n330, Q => 
                           REGISTERS_28_14_port, QN => n_5358);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => n324, Q => 
                           REGISTERS_28_13_port, QN => n_5359);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => n321, Q => 
                           REGISTERS_28_12_port, QN => n_5360);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => n317, Q => 
                           REGISTERS_28_11_port, QN => n_5361);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => n314, Q => 
                           REGISTERS_28_10_port, QN => n_5362);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => n311, Q => 
                           REGISTERS_28_9_port, QN => n_5363);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => n308, Q => 
                           REGISTERS_28_8_port, QN => n_5364);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => n305, Q => 
                           REGISTERS_28_7_port, QN => n_5365);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => n302, Q => 
                           REGISTERS_28_6_port, QN => n_5366);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => n299, Q => 
                           REGISTERS_28_5_port, QN => n_5367);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => n296, Q => 
                           REGISTERS_28_4_port, QN => n_5368);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => n293, Q => 
                           REGISTERS_28_3_port, QN => n_5369);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => n364, Q => 
                           REGISTERS_28_2_port, QN => n_5370);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => n290, Q => 
                           REGISTERS_28_1_port, QN => n_5371);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => n370, Q => 
                           REGISTERS_28_0_port, QN => n_5372);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => n373, Q => 
                           REGISTERS_29_31_port, QN => n_5373);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => n376, Q => 
                           REGISTERS_29_30_port, QN => n_5374);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => n379, Q => 
                           REGISTERS_29_29_port, QN => n_5375);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => n382, Q => 
                           REGISTERS_29_28_port, QN => n_5376);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => n385_port, Q 
                           => REGISTERS_29_27_port, QN => n_5377);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => n367, Q => 
                           REGISTERS_29_26_port, QN => n_5378);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => n354, Q => 
                           REGISTERS_29_25_port, QN => n_5379);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => n357, Q => 
                           REGISTERS_29_24_port, QN => n_5380);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => n345, Q => 
                           REGISTERS_29_23_port, QN => n_5381);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => n348, Q => 
                           REGISTERS_29_22_port, QN => n_5382);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => n351, Q => 
                           REGISTERS_29_21_port, QN => n_5383);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => n333, Q => 
                           REGISTERS_29_20_port, QN => n_5384);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => n336, Q => 
                           REGISTERS_29_19_port, QN => n_5385);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => n339, Q => 
                           REGISTERS_29_18_port, QN => n_5386);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => n361, Q => 
                           REGISTERS_29_17_port, QN => n_5387);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => n342, Q => 
                           REGISTERS_29_16_port, QN => n_5388);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => n327, Q => 
                           REGISTERS_29_15_port, QN => n_5389);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => n330, Q => 
                           REGISTERS_29_14_port, QN => n_5390);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => n324, Q => 
                           REGISTERS_29_13_port, QN => n_5391);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => n321, Q => 
                           REGISTERS_29_12_port, QN => n_5392);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => n318, Q => 
                           REGISTERS_29_11_port, QN => n_5393);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => n314, Q => 
                           REGISTERS_29_10_port, QN => n_5394);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => n311, Q => 
                           REGISTERS_29_9_port, QN => n_5395);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => n308, Q => 
                           REGISTERS_29_8_port, QN => n_5396);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => n305, Q => 
                           REGISTERS_29_7_port, QN => n_5397);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => n302, Q => 
                           REGISTERS_29_6_port, QN => n_5398);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => n299, Q => 
                           REGISTERS_29_5_port, QN => n_5399);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => n296, Q => 
                           REGISTERS_29_4_port, QN => n_5400);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => n293, Q => 
                           REGISTERS_29_3_port, QN => n_5401);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => n364, Q => 
                           REGISTERS_29_2_port, QN => n_5402);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => n290, Q => 
                           REGISTERS_29_1_port, QN => n_5403);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => n370, Q => 
                           REGISTERS_29_0_port, QN => n_5404);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => n373, Q => 
                           REGISTERS_30_31_port, QN => n_5405);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => n376, Q => 
                           REGISTERS_30_30_port, QN => n_5406);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => n379, Q => 
                           REGISTERS_30_29_port, QN => n_5407);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => n382, Q => 
                           REGISTERS_30_28_port, QN => n_5408);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => n385_port, Q 
                           => REGISTERS_30_27_port, QN => n_5409);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => n367, Q => 
                           REGISTERS_30_26_port, QN => n_5410);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => n354, Q => 
                           REGISTERS_30_25_port, QN => n_5411);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => n358, Q => 
                           REGISTERS_30_24_port, QN => n_5412);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => n345, Q => 
                           REGISTERS_30_23_port, QN => n_5413);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => n348, Q => 
                           REGISTERS_30_22_port, QN => n_5414);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => n351, Q => 
                           REGISTERS_30_21_port, QN => n_5415);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => n333, Q => 
                           REGISTERS_30_20_port, QN => n_5416);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => n336, Q => 
                           REGISTERS_30_19_port, QN => n_5417);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => n339, Q => 
                           REGISTERS_30_18_port, QN => n_5418);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => n361, Q => 
                           REGISTERS_30_17_port, QN => n_5419);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => n342, Q => 
                           REGISTERS_30_16_port, QN => n_5420);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => n327, Q => 
                           REGISTERS_30_15_port, QN => n_5421);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => n330, Q => 
                           REGISTERS_30_14_port, QN => n_5422);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => n324, Q => 
                           REGISTERS_30_13_port, QN => n_5423);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => n321, Q => 
                           REGISTERS_30_12_port, QN => n_5424);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => n318, Q => 
                           REGISTERS_30_11_port, QN => n_5425);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => n315, Q => 
                           REGISTERS_30_10_port, QN => n_5426);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => n311, Q => 
                           REGISTERS_30_9_port, QN => n_5427);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => n308, Q => 
                           REGISTERS_30_8_port, QN => n_5428);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => n305, Q => 
                           REGISTERS_30_7_port, QN => n_5429);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => n302, Q => 
                           REGISTERS_30_6_port, QN => n_5430);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => n299, Q => 
                           REGISTERS_30_5_port, QN => n_5431);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => n296, Q => 
                           REGISTERS_30_4_port, QN => n_5432);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => n293, Q => 
                           REGISTERS_30_3_port, QN => n_5433);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => n364, Q => 
                           REGISTERS_30_2_port, QN => n_5434);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => n290, Q => 
                           REGISTERS_30_1_port, QN => n_5435);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => n370, Q => 
                           REGISTERS_30_0_port, QN => n_5436);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => n373, Q => 
                           REGISTERS_31_31_port, QN => n_5437);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => n376, Q => 
                           REGISTERS_31_30_port, QN => n_5438);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => n379, Q => 
                           REGISTERS_31_29_port, QN => n_5439);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => n382, Q => 
                           REGISTERS_31_28_port, QN => n_5440);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => n385_port, Q 
                           => REGISTERS_31_27_port, QN => n_5441);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => n367, Q => 
                           REGISTERS_31_26_port, QN => n_5442);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => n355, Q => 
                           REGISTERS_31_25_port, QN => n_5443);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => n358, Q => 
                           REGISTERS_31_24_port, QN => n_5444);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => n345, Q => 
                           REGISTERS_31_23_port, QN => n_5445);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => n348, Q => 
                           REGISTERS_31_22_port, QN => n_5446);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => n352, Q => 
                           REGISTERS_31_21_port, QN => n_5447);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => n333, Q => 
                           REGISTERS_31_20_port, QN => n_5448);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => n336, Q => 
                           REGISTERS_31_19_port, QN => n_5449);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => n339, Q => 
                           REGISTERS_31_18_port, QN => n_5450);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => n361, Q => 
                           REGISTERS_31_17_port, QN => n_5451);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => n342, Q => 
                           REGISTERS_31_16_port, QN => n_5452);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => n327, Q => 
                           REGISTERS_31_15_port, QN => n_5453);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => n330, Q => 
                           REGISTERS_31_14_port, QN => n_5454);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => n324, Q => 
                           REGISTERS_31_13_port, QN => n_5455);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => n321, Q => 
                           REGISTERS_31_12_port, QN => n_5456);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => n318, Q => 
                           REGISTERS_31_11_port, QN => n_5457);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => n315, Q => 
                           REGISTERS_31_10_port, QN => n_5458);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => n312, Q => 
                           REGISTERS_31_9_port, QN => n_5459);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => n308, Q => 
                           REGISTERS_31_8_port, QN => n_5460);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => n305, Q => 
                           REGISTERS_31_7_port, QN => n_5461);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => n302, Q => 
                           REGISTERS_31_6_port, QN => n_5462);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => n299, Q => 
                           REGISTERS_31_5_port, QN => n_5463);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => n296, Q => 
                           REGISTERS_31_4_port, QN => n_5464);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => n293, Q => 
                           REGISTERS_31_3_port, QN => n_5465);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => n364, Q => 
                           REGISTERS_31_2_port, QN => n_5466);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => n290, Q => 
                           REGISTERS_31_1_port, QN => n_5467);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => n370, Q => 
                           REGISTERS_31_0_port, QN => n_5468);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => n370, Q => OUT1(31), QN
                           => n_5469);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => n373, Q => OUT1(30), QN
                           => n_5470);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => n376, Q => OUT1(29), QN
                           => n_5471);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => n379, Q => OUT1(28), QN
                           => n_5472);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => n382, Q => OUT1(27), QN
                           => n_5473);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => n364, Q => OUT1(26), QN
                           => n_5474);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => n352, Q => OUT1(25), QN
                           => n_5475);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => n355, Q => OUT1(24), QN
                           => n_5476);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => n342, Q => OUT1(23), QN
                           => n_5477);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => n346, Q => OUT1(22), QN
                           => n_5478);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => n349, Q => OUT1(21), QN
                           => n_5479);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => n330, Q => OUT1(20), QN
                           => n_5480);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => n333, Q => OUT1(19), QN
                           => n_5481);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => n336, Q => OUT1(18), QN
                           => n_5482);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => n358, Q => OUT1(17), QN
                           => n_5483);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => n339, Q => OUT1(16), QN
                           => n_5484);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => n324, Q => OUT1(15), QN
                           => n_5485);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => n327, Q => OUT1(14), QN
                           => n_5486);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => n321, Q => OUT1(13), QN
                           => n_5487);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => n318, Q => OUT1(12), QN
                           => n_5488);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => n315, Q => OUT1(11), QN
                           => n_5489);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => n312, Q => OUT1(10), QN
                           => n_5490);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => n309, Q => OUT1(9), QN 
                           => n_5491);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => n306, Q => OUT1(8), QN 
                           => n_5492);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => n302, Q => OUT1(7), QN 
                           => n_5493);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => n299, Q => OUT1(6), QN 
                           => n_5494);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => n296, Q => OUT1(5), QN 
                           => n_5495);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => n293, Q => OUT1(4), QN 
                           => n_5496);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => n290, Q => OUT1(3), QN 
                           => n_5497);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => n361, Q => OUT1(2), QN 
                           => n_5498);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => n287, Q => OUT1(1), QN 
                           => n_5499);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => n367, Q => OUT1(0), QN 
                           => n_5500);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => n370, Q => OUT2(31), QN
                           => n_5501);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => n373, Q => OUT2(30), QN
                           => n_5502);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => n376, Q => OUT2(29), QN
                           => n_5503);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => n379, Q => OUT2(28), QN
                           => n_5504);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => n382, Q => OUT2(27), QN
                           => n_5505);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => n287, Q => OUT2(26), QN
                           => n_5506);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => n287, Q => OUT2(25), QN
                           => n_5507);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => n355, Q => OUT2(24), QN
                           => n_5508);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => n287, Q => OUT2(23), QN
                           => n_5509);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => n345, Q => OUT2(22), QN
                           => n_5510);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => n349, Q => OUT2(21), QN
                           => n_5511);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => n287, Q => OUT2(20), QN
                           => n_5512);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => n333, Q => OUT2(19), QN
                           => n_5513);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => n336, Q => OUT2(18), QN
                           => n_5514);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => n358, Q => OUT2(17), QN
                           => n_5515);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => n339, Q => OUT2(16), QN
                           => n_5516);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => n324, Q => OUT2(15), QN
                           => n_5517);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => n327, Q => OUT2(14), QN
                           => n_5518);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => n321, Q => OUT2(13), QN
                           => n_5519);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => n318, Q => OUT2(12), QN
                           => n_5520);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => n315, Q => OUT2(11), QN
                           => n_5521);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => n312, Q => OUT2(10), QN
                           => n_5522);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => n309, Q => OUT2(9), QN 
                           => n_5523);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => n305, Q => OUT2(8), QN 
                           => n_5524);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => n302, Q => OUT2(7), QN 
                           => n_5525);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => n299, Q => OUT2(6), QN 
                           => n_5526);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => n296, Q => OUT2(5), QN 
                           => n_5527);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => n293, Q => OUT2(4), QN 
                           => n_5528);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => n290, Q => OUT2(3), QN 
                           => n_5529);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => n361, Q => OUT2(2), QN 
                           => n_5530);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => n287, Q => OUT2(1), QN 
                           => n_5531);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => n367, Q => OUT2(0), QN 
                           => n_5532);
   U3 : INV_X1 port map( A => n2869, ZN => n1);
   U4 : INV_X2 port map( A => n1, ZN => n2);
   U5 : INV_X1 port map( A => n2870, ZN => n3);
   U6 : INV_X2 port map( A => n3, ZN => n4);
   U7 : INV_X1 port map( A => n2871, ZN => n5);
   U8 : INV_X2 port map( A => n5, ZN => n6);
   U9 : INV_X1 port map( A => n2872, ZN => n7);
   U10 : INV_X2 port map( A => n7, ZN => n8);
   U11 : INV_X1 port map( A => n2874, ZN => n9);
   U12 : INV_X2 port map( A => n9, ZN => n10);
   U13 : INV_X1 port map( A => n2875, ZN => n11);
   U14 : INV_X2 port map( A => n11, ZN => n12);
   U15 : INV_X1 port map( A => n2876, ZN => n13);
   U16 : INV_X2 port map( A => n13, ZN => n14);
   U17 : INV_X1 port map( A => n2877, ZN => n15);
   U18 : INV_X2 port map( A => n15, ZN => n16);
   U19 : INV_X1 port map( A => n2878, ZN => n17);
   U20 : INV_X2 port map( A => n17, ZN => n18);
   U21 : INV_X1 port map( A => n2879, ZN => n19);
   U22 : INV_X2 port map( A => n19, ZN => n20);
   U23 : INV_X1 port map( A => n2880, ZN => n21);
   U24 : INV_X2 port map( A => n21, ZN => n22);
   U25 : INV_X1 port map( A => n2881, ZN => n23);
   U26 : INV_X2 port map( A => n23, ZN => n24);
   U27 : INV_X1 port map( A => n2886, ZN => n25);
   U28 : INV_X2 port map( A => n25, ZN => n26);
   U29 : INV_X1 port map( A => n2887, ZN => n27);
   U30 : INV_X2 port map( A => n27, ZN => n28);
   U31 : INV_X1 port map( A => n2888, ZN => n29);
   U32 : INV_X2 port map( A => n29, ZN => n30);
   U33 : INV_X1 port map( A => n2889, ZN => n31_port);
   U34 : INV_X2 port map( A => n31_port, ZN => n32_port);
   U35 : INV_X1 port map( A => n2890, ZN => n33_port);
   U36 : INV_X2 port map( A => n33_port, ZN => n34_port);
   U37 : INV_X1 port map( A => n2891, ZN => n35_port);
   U38 : INV_X2 port map( A => n35_port, ZN => n36_port);
   U39 : INV_X1 port map( A => n2892, ZN => n37_port);
   U40 : INV_X2 port map( A => n37_port, ZN => n38_port);
   U41 : INV_X1 port map( A => n2867, ZN => n39_port);
   U42 : INV_X2 port map( A => n39_port, ZN => n40_port);
   U43 : INV_X1 port map( A => n2868, ZN => n41_port);
   U44 : INV_X2 port map( A => n41_port, ZN => n42_port);
   U45 : INV_X1 port map( A => n2865, ZN => n43_port);
   U46 : INV_X2 port map( A => n43_port, ZN => n44_port);
   U47 : INV_X1 port map( A => n2866, ZN => n45_port);
   U48 : INV_X2 port map( A => n45_port, ZN => n46_port);
   U49 : INV_X1 port map( A => n2858, ZN => n47_port);
   U50 : INV_X2 port map( A => n47_port, ZN => n48_port);
   U51 : INV_X1 port map( A => n2863, ZN => n49_port);
   U52 : INV_X2 port map( A => n49_port, ZN => n50_port);
   U53 : INV_X1 port map( A => n2854, ZN => n51_port);
   U54 : INV_X2 port map( A => n51_port, ZN => n52_port);
   U55 : INV_X1 port map( A => n2856, ZN => n53_port);
   U56 : INV_X2 port map( A => n53_port, ZN => n54_port);
   U57 : INV_X1 port map( A => n2850, ZN => n55_port);
   U58 : INV_X2 port map( A => n55_port, ZN => n56_port);
   U59 : INV_X1 port map( A => n2852, ZN => n57_port);
   U60 : INV_X2 port map( A => n57_port, ZN => n58_port);
   U61 : INV_X1 port map( A => n2846, ZN => n59_port);
   U62 : INV_X2 port map( A => n59_port, ZN => n60_port);
   U63 : INV_X1 port map( A => n2848, ZN => n61_port);
   U64 : INV_X2 port map( A => n61_port, ZN => n62_port);
   U65 : INV_X1 port map( A => n2812, ZN => n63);
   U66 : INV_X2 port map( A => n63, ZN => n64);
   U67 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1087);
   U68 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n2803);
   U69 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => n1091, ZN => n1089);
   U70 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => n2807, ZN => n2805);
   U71 : NOR2_X4 port map( A1 => n1091, A2 => ADD_RD1(4), ZN => n1083);
   U72 : NOR2_X4 port map( A1 => n2807, A2 => ADD_RD2(4), ZN => n2799);
   U73 : NOR2_X4 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1085);
   U74 : NOR2_X4 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n2801);
   U75 : BUF_X1 port map( A => n283, Z => n400_port);
   U76 : BUF_X1 port map( A => n283, Z => n399_port);
   U77 : BUF_X1 port map( A => n283, Z => n398_port);
   U78 : BUF_X1 port map( A => n282, Z => n397_port);
   U79 : BUF_X1 port map( A => n282, Z => n396_port);
   U80 : BUF_X1 port map( A => n280, Z => n390_port);
   U81 : BUF_X1 port map( A => n281, Z => n394_port);
   U82 : BUF_X1 port map( A => n282, Z => n395_port);
   U83 : BUF_X1 port map( A => n281, Z => n392_port);
   U84 : BUF_X1 port map( A => n281, Z => n393_port);
   U85 : BUF_X1 port map( A => n280, Z => n391_port);
   U86 : BUF_X1 port map( A => n280, Z => n389_port);
   U87 : BUF_X1 port map( A => n279, Z => n386_port);
   U88 : BUF_X1 port map( A => n279, Z => n387_port);
   U89 : BUF_X1 port map( A => n279, Z => n388_port);
   U90 : BUF_X1 port map( A => n284, Z => n401_port);
   U91 : BUF_X1 port map( A => n284, Z => n402_port);
   U92 : BUF_X1 port map( A => n2793, Z => n260);
   U93 : BUF_X1 port map( A => n2792, Z => n247);
   U94 : BUF_X1 port map( A => n2791, Z => n234);
   U95 : BUF_X1 port map( A => n2790, Z => n221);
   U96 : BUF_X1 port map( A => n1077, Z => n156);
   U97 : BUF_X1 port map( A => n1076, Z => n143);
   U98 : BUF_X1 port map( A => n1075, Z => n130);
   U99 : BUF_X1 port map( A => n1074, Z => n117_port);
   U100 : BUF_X1 port map( A => n2793, Z => n261);
   U101 : BUF_X1 port map( A => n2792, Z => n248);
   U102 : BUF_X1 port map( A => n2791, Z => n235);
   U103 : BUF_X1 port map( A => n2790, Z => n222);
   U104 : BUF_X1 port map( A => n1077, Z => n157);
   U105 : BUF_X1 port map( A => n1076, Z => n144);
   U106 : BUF_X1 port map( A => n1075, Z => n131);
   U107 : BUF_X1 port map( A => n1074, Z => n118_port);
   U108 : BUF_X1 port map( A => n285, Z => n283);
   U109 : BUF_X1 port map( A => n285, Z => n282);
   U110 : BUF_X1 port map( A => n286, Z => n281);
   U111 : BUF_X1 port map( A => n286, Z => n280);
   U112 : BUF_X1 port map( A => n286, Z => n279);
   U113 : BUF_X1 port map( A => n285, Z => n284);
   U114 : INV_X1 port map( A => RESET, ZN => n278);
   U115 : BUF_X1 port map( A => CLK, Z => n285);
   U116 : BUF_X1 port map( A => CLK, Z => n286);
   U117 : BUF_X1 port map( A => n2786, Z => n169);
   U118 : BUF_X1 port map( A => n2789, Z => n208);
   U119 : BUF_X1 port map( A => n2788, Z => n195);
   U120 : BUF_X1 port map( A => n2787, Z => n182);
   U121 : BUF_X1 port map( A => n1070, Z => n65);
   U122 : BUF_X1 port map( A => n1073, Z => n104_port);
   U123 : BUF_X1 port map( A => n1072, Z => n91);
   U124 : BUF_X1 port map( A => n1071, Z => n78);
   U125 : BUF_X1 port map( A => n2786, Z => n170);
   U126 : BUF_X1 port map( A => n2789, Z => n209);
   U127 : BUF_X1 port map( A => n2788, Z => n196);
   U128 : BUF_X1 port map( A => n2787, Z => n183);
   U129 : BUF_X1 port map( A => n1070, Z => n66);
   U130 : BUF_X1 port map( A => n1073, Z => n105_port);
   U131 : BUF_X1 port map( A => n1072, Z => n92);
   U132 : BUF_X1 port map( A => n1071, Z => n79);
   U133 : INV_X1 port map( A => ADD_RD2(0), ZN => n2810);
   U134 : INV_X1 port map( A => ADD_RD1(0), ZN => n1094);
   U135 : INV_X1 port map( A => ADD_RD2(2), ZN => n2808);
   U136 : INV_X1 port map( A => ADD_RD2(3), ZN => n2807);
   U137 : INV_X1 port map( A => ADD_RD2(1), ZN => n2809);
   U138 : INV_X1 port map( A => ADD_RD1(2), ZN => n1092);
   U139 : INV_X1 port map( A => ADD_RD1(3), ZN => n1091);
   U140 : INV_X1 port map( A => ADD_RD1(1), ZN => n1093);
   U141 : CLKBUF_X1 port map( A => n65, Z => n67);
   U142 : CLKBUF_X1 port map( A => n65, Z => n68);
   U143 : CLKBUF_X1 port map( A => n65, Z => n69);
   U144 : CLKBUF_X1 port map( A => n65, Z => n70);
   U145 : CLKBUF_X1 port map( A => n65, Z => n71);
   U146 : CLKBUF_X1 port map( A => n65, Z => n72);
   U147 : CLKBUF_X1 port map( A => n66, Z => n73);
   U148 : CLKBUF_X1 port map( A => n66, Z => n74);
   U149 : CLKBUF_X1 port map( A => n66, Z => n75);
   U150 : CLKBUF_X1 port map( A => n66, Z => n76);
   U151 : CLKBUF_X1 port map( A => n66, Z => n77);
   U152 : CLKBUF_X1 port map( A => n78, Z => n80);
   U153 : CLKBUF_X1 port map( A => n78, Z => n81);
   U154 : CLKBUF_X1 port map( A => n78, Z => n82);
   U155 : CLKBUF_X1 port map( A => n78, Z => n83);
   U156 : CLKBUF_X1 port map( A => n78, Z => n84);
   U157 : CLKBUF_X1 port map( A => n78, Z => n85);
   U158 : CLKBUF_X1 port map( A => n79, Z => n86);
   U159 : CLKBUF_X1 port map( A => n79, Z => n87);
   U160 : CLKBUF_X1 port map( A => n79, Z => n88);
   U161 : CLKBUF_X1 port map( A => n79, Z => n89);
   U162 : CLKBUF_X1 port map( A => n79, Z => n90);
   U163 : CLKBUF_X1 port map( A => n91, Z => n93);
   U164 : CLKBUF_X1 port map( A => n91, Z => n94);
   U165 : CLKBUF_X1 port map( A => n91, Z => n95);
   U166 : CLKBUF_X1 port map( A => n91, Z => n96_port);
   U167 : CLKBUF_X1 port map( A => n91, Z => n97_port);
   U168 : CLKBUF_X1 port map( A => n91, Z => n98_port);
   U169 : CLKBUF_X1 port map( A => n92, Z => n99_port);
   U170 : CLKBUF_X1 port map( A => n92, Z => n100_port);
   U171 : CLKBUF_X1 port map( A => n92, Z => n101_port);
   U172 : CLKBUF_X1 port map( A => n92, Z => n102_port);
   U173 : CLKBUF_X1 port map( A => n92, Z => n103_port);
   U174 : CLKBUF_X1 port map( A => n104_port, Z => n106_port);
   U175 : CLKBUF_X1 port map( A => n104_port, Z => n107_port);
   U176 : CLKBUF_X1 port map( A => n104_port, Z => n108_port);
   U177 : CLKBUF_X1 port map( A => n104_port, Z => n109_port);
   U178 : CLKBUF_X1 port map( A => n104_port, Z => n110_port);
   U179 : CLKBUF_X1 port map( A => n104_port, Z => n111_port);
   U180 : CLKBUF_X1 port map( A => n105_port, Z => n112_port);
   U181 : CLKBUF_X1 port map( A => n105_port, Z => n113_port);
   U182 : CLKBUF_X1 port map( A => n105_port, Z => n114_port);
   U183 : CLKBUF_X1 port map( A => n105_port, Z => n115_port);
   U184 : CLKBUF_X1 port map( A => n105_port, Z => n116_port);
   U185 : CLKBUF_X1 port map( A => n117_port, Z => n119_port);
   U186 : CLKBUF_X1 port map( A => n117_port, Z => n120_port);
   U187 : CLKBUF_X1 port map( A => n117_port, Z => n121_port);
   U188 : CLKBUF_X1 port map( A => n117_port, Z => n122_port);
   U189 : CLKBUF_X1 port map( A => n117_port, Z => n123_port);
   U190 : CLKBUF_X1 port map( A => n117_port, Z => n124_port);
   U191 : CLKBUF_X1 port map( A => n118_port, Z => n125_port);
   U192 : CLKBUF_X1 port map( A => n118_port, Z => n126_port);
   U193 : CLKBUF_X1 port map( A => n118_port, Z => n127_port);
   U194 : CLKBUF_X1 port map( A => n118_port, Z => n128);
   U195 : CLKBUF_X1 port map( A => n118_port, Z => n129);
   U196 : CLKBUF_X1 port map( A => n130, Z => n132);
   U197 : CLKBUF_X1 port map( A => n130, Z => n133);
   U198 : CLKBUF_X1 port map( A => n130, Z => n134);
   U199 : CLKBUF_X1 port map( A => n130, Z => n135);
   U200 : CLKBUF_X1 port map( A => n130, Z => n136);
   U201 : CLKBUF_X1 port map( A => n130, Z => n137);
   U202 : CLKBUF_X1 port map( A => n131, Z => n138);
   U203 : CLKBUF_X1 port map( A => n131, Z => n139);
   U204 : CLKBUF_X1 port map( A => n131, Z => n140);
   U205 : CLKBUF_X1 port map( A => n131, Z => n141);
   U206 : CLKBUF_X1 port map( A => n131, Z => n142);
   U207 : CLKBUF_X1 port map( A => n143, Z => n145);
   U208 : CLKBUF_X1 port map( A => n143, Z => n146);
   U209 : CLKBUF_X1 port map( A => n143, Z => n147);
   U210 : CLKBUF_X1 port map( A => n143, Z => n148);
   U211 : CLKBUF_X1 port map( A => n143, Z => n149);
   U212 : CLKBUF_X1 port map( A => n143, Z => n150);
   U213 : CLKBUF_X1 port map( A => n144, Z => n151);
   U214 : CLKBUF_X1 port map( A => n144, Z => n152);
   U215 : CLKBUF_X1 port map( A => n144, Z => n153);
   U216 : CLKBUF_X1 port map( A => n144, Z => n154);
   U217 : CLKBUF_X1 port map( A => n144, Z => n155);
   U218 : CLKBUF_X1 port map( A => n156, Z => n158);
   U219 : CLKBUF_X1 port map( A => n156, Z => n159);
   U220 : CLKBUF_X1 port map( A => n156, Z => n160);
   U221 : CLKBUF_X1 port map( A => n156, Z => n161);
   U222 : CLKBUF_X1 port map( A => n156, Z => n162);
   U223 : CLKBUF_X1 port map( A => n156, Z => n163);
   U224 : CLKBUF_X1 port map( A => n157, Z => n164);
   U225 : CLKBUF_X1 port map( A => n157, Z => n165);
   U226 : CLKBUF_X1 port map( A => n157, Z => n166);
   U227 : CLKBUF_X1 port map( A => n157, Z => n167);
   U228 : CLKBUF_X1 port map( A => n157, Z => n168);
   U229 : CLKBUF_X1 port map( A => n169, Z => n171);
   U230 : CLKBUF_X1 port map( A => n169, Z => n172);
   U231 : CLKBUF_X1 port map( A => n169, Z => n173);
   U232 : CLKBUF_X1 port map( A => n169, Z => n174);
   U233 : CLKBUF_X1 port map( A => n169, Z => n175);
   U234 : CLKBUF_X1 port map( A => n169, Z => n176);
   U235 : CLKBUF_X1 port map( A => n170, Z => n177);
   U236 : CLKBUF_X1 port map( A => n170, Z => n178);
   U237 : CLKBUF_X1 port map( A => n170, Z => n179);
   U238 : CLKBUF_X1 port map( A => n170, Z => n180);
   U239 : CLKBUF_X1 port map( A => n170, Z => n181);
   U240 : CLKBUF_X1 port map( A => n182, Z => n184);
   U241 : CLKBUF_X1 port map( A => n182, Z => n185);
   U242 : CLKBUF_X1 port map( A => n182, Z => n186);
   U243 : CLKBUF_X1 port map( A => n182, Z => n187);
   U244 : CLKBUF_X1 port map( A => n182, Z => n188);
   U245 : CLKBUF_X1 port map( A => n182, Z => n189);
   U246 : CLKBUF_X1 port map( A => n183, Z => n190);
   U247 : CLKBUF_X1 port map( A => n183, Z => n191);
   U248 : CLKBUF_X1 port map( A => n183, Z => n192);
   U249 : CLKBUF_X1 port map( A => n183, Z => n193);
   U250 : CLKBUF_X1 port map( A => n183, Z => n194);
   U251 : CLKBUF_X1 port map( A => n195, Z => n197);
   U252 : CLKBUF_X1 port map( A => n195, Z => n198);
   U253 : CLKBUF_X1 port map( A => n195, Z => n199);
   U254 : CLKBUF_X1 port map( A => n195, Z => n200);
   U255 : CLKBUF_X1 port map( A => n195, Z => n201);
   U256 : CLKBUF_X1 port map( A => n195, Z => n202);
   U257 : CLKBUF_X1 port map( A => n196, Z => n203);
   U258 : CLKBUF_X1 port map( A => n196, Z => n204);
   U259 : CLKBUF_X1 port map( A => n196, Z => n205);
   U260 : CLKBUF_X1 port map( A => n196, Z => n206);
   U261 : CLKBUF_X1 port map( A => n196, Z => n207);
   U262 : CLKBUF_X1 port map( A => n208, Z => n210);
   U263 : CLKBUF_X1 port map( A => n208, Z => n211);
   U264 : CLKBUF_X1 port map( A => n208, Z => n212);
   U265 : CLKBUF_X1 port map( A => n208, Z => n213);
   U266 : CLKBUF_X1 port map( A => n208, Z => n214);
   U267 : CLKBUF_X1 port map( A => n208, Z => n215);
   U268 : CLKBUF_X1 port map( A => n209, Z => n216);
   U269 : CLKBUF_X1 port map( A => n209, Z => n217);
   U270 : CLKBUF_X1 port map( A => n209, Z => n218);
   U271 : CLKBUF_X1 port map( A => n209, Z => n219);
   U272 : CLKBUF_X1 port map( A => n209, Z => n220);
   U273 : CLKBUF_X1 port map( A => n221, Z => n223);
   U274 : CLKBUF_X1 port map( A => n221, Z => n224);
   U275 : CLKBUF_X1 port map( A => n221, Z => n225);
   U276 : CLKBUF_X1 port map( A => n221, Z => n226);
   U277 : CLKBUF_X1 port map( A => n221, Z => n227);
   U278 : CLKBUF_X1 port map( A => n221, Z => n228);
   U279 : CLKBUF_X1 port map( A => n222, Z => n229);
   U280 : CLKBUF_X1 port map( A => n222, Z => n230);
   U281 : CLKBUF_X1 port map( A => n222, Z => n231);
   U282 : CLKBUF_X1 port map( A => n222, Z => n232);
   U283 : CLKBUF_X1 port map( A => n222, Z => n233);
   U284 : CLKBUF_X1 port map( A => n234, Z => n236);
   U285 : CLKBUF_X1 port map( A => n234, Z => n237);
   U286 : CLKBUF_X1 port map( A => n234, Z => n238);
   U287 : CLKBUF_X1 port map( A => n234, Z => n239);
   U288 : CLKBUF_X1 port map( A => n234, Z => n240);
   U289 : CLKBUF_X1 port map( A => n234, Z => n241);
   U290 : CLKBUF_X1 port map( A => n235, Z => n242);
   U291 : CLKBUF_X1 port map( A => n235, Z => n243);
   U292 : CLKBUF_X1 port map( A => n235, Z => n244);
   U293 : CLKBUF_X1 port map( A => n235, Z => n245);
   U294 : CLKBUF_X1 port map( A => n235, Z => n246);
   U295 : CLKBUF_X1 port map( A => n247, Z => n249);
   U296 : CLKBUF_X1 port map( A => n247, Z => n250);
   U297 : CLKBUF_X1 port map( A => n247, Z => n251);
   U298 : CLKBUF_X1 port map( A => n247, Z => n252);
   U299 : CLKBUF_X1 port map( A => n247, Z => n253);
   U300 : CLKBUF_X1 port map( A => n247, Z => n254);
   U301 : CLKBUF_X1 port map( A => n248, Z => n255);
   U302 : CLKBUF_X1 port map( A => n248, Z => n256);
   U303 : CLKBUF_X1 port map( A => n248, Z => n257);
   U304 : CLKBUF_X1 port map( A => n248, Z => n258);
   U305 : CLKBUF_X1 port map( A => n248, Z => n259);
   U306 : CLKBUF_X1 port map( A => n260, Z => n262);
   U307 : CLKBUF_X1 port map( A => n260, Z => n263);
   U308 : CLKBUF_X1 port map( A => n260, Z => n264);
   U309 : CLKBUF_X1 port map( A => n260, Z => n265);
   U310 : CLKBUF_X1 port map( A => n260, Z => n266);
   U311 : CLKBUF_X1 port map( A => n260, Z => n267);
   U312 : CLKBUF_X1 port map( A => n261, Z => n268);
   U313 : CLKBUF_X1 port map( A => n261, Z => n269);
   U314 : CLKBUF_X1 port map( A => n261, Z => n270);
   U315 : CLKBUF_X1 port map( A => n261, Z => n271);
   U316 : CLKBUF_X1 port map( A => n261, Z => n272);
   U317 : CLKBUF_X1 port map( A => n278, Z => n273);
   U318 : CLKBUF_X1 port map( A => n278, Z => n274);
   U319 : CLKBUF_X1 port map( A => n278, Z => n275);
   U320 : CLKBUF_X1 port map( A => n278, Z => n276);
   U321 : CLKBUF_X1 port map( A => n278, Z => n277);
   U322 : CLKBUF_X1 port map( A => n402_port, Z => n287);
   U323 : CLKBUF_X1 port map( A => n402_port, Z => n288);
   U324 : CLKBUF_X1 port map( A => n402_port, Z => n289);
   U325 : CLKBUF_X1 port map( A => n401_port, Z => n290);
   U326 : CLKBUF_X1 port map( A => n401_port, Z => n291);
   U327 : CLKBUF_X1 port map( A => n401_port, Z => n292);
   U328 : CLKBUF_X1 port map( A => n401_port, Z => n293);
   U329 : CLKBUF_X1 port map( A => n401_port, Z => n294);
   U330 : CLKBUF_X1 port map( A => n401_port, Z => n295);
   U331 : CLKBUF_X1 port map( A => n400_port, Z => n296);
   U332 : CLKBUF_X1 port map( A => n400_port, Z => n297);
   U333 : CLKBUF_X1 port map( A => n400_port, Z => n298);
   U334 : CLKBUF_X1 port map( A => n400_port, Z => n299);
   U335 : CLKBUF_X1 port map( A => n400_port, Z => n300);
   U336 : CLKBUF_X1 port map( A => n400_port, Z => n301);
   U337 : CLKBUF_X1 port map( A => n399_port, Z => n302);
   U338 : CLKBUF_X1 port map( A => n399_port, Z => n303);
   U339 : CLKBUF_X1 port map( A => n399_port, Z => n304);
   U340 : CLKBUF_X1 port map( A => n399_port, Z => n305);
   U341 : CLKBUF_X1 port map( A => n399_port, Z => n306);
   U342 : CLKBUF_X1 port map( A => n399_port, Z => n307);
   U343 : CLKBUF_X1 port map( A => n398_port, Z => n308);
   U344 : CLKBUF_X1 port map( A => n398_port, Z => n309);
   U345 : CLKBUF_X1 port map( A => n398_port, Z => n310);
   U346 : CLKBUF_X1 port map( A => n398_port, Z => n311);
   U347 : CLKBUF_X1 port map( A => n398_port, Z => n312);
   U348 : CLKBUF_X1 port map( A => n398_port, Z => n313);
   U349 : CLKBUF_X1 port map( A => n397_port, Z => n314);
   U350 : CLKBUF_X1 port map( A => n397_port, Z => n315);
   U351 : CLKBUF_X1 port map( A => n397_port, Z => n316);
   U352 : CLKBUF_X1 port map( A => n397_port, Z => n317);
   U353 : CLKBUF_X1 port map( A => n397_port, Z => n318);
   U354 : CLKBUF_X1 port map( A => n397_port, Z => n319);
   U355 : CLKBUF_X1 port map( A => n396_port, Z => n320);
   U356 : CLKBUF_X1 port map( A => n396_port, Z => n321);
   U357 : CLKBUF_X1 port map( A => n396_port, Z => n322);
   U358 : CLKBUF_X1 port map( A => n396_port, Z => n323);
   U359 : CLKBUF_X1 port map( A => n396_port, Z => n324);
   U360 : CLKBUF_X1 port map( A => n396_port, Z => n325);
   U361 : CLKBUF_X1 port map( A => n395_port, Z => n326);
   U362 : CLKBUF_X1 port map( A => n395_port, Z => n327);
   U363 : CLKBUF_X1 port map( A => n395_port, Z => n328);
   U364 : CLKBUF_X1 port map( A => n395_port, Z => n329);
   U365 : CLKBUF_X1 port map( A => n395_port, Z => n330);
   U366 : CLKBUF_X1 port map( A => n395_port, Z => n331);
   U367 : CLKBUF_X1 port map( A => n394_port, Z => n332);
   U368 : CLKBUF_X1 port map( A => n394_port, Z => n333);
   U369 : CLKBUF_X1 port map( A => n394_port, Z => n334);
   U370 : CLKBUF_X1 port map( A => n394_port, Z => n335);
   U371 : CLKBUF_X1 port map( A => n394_port, Z => n336);
   U372 : CLKBUF_X1 port map( A => n394_port, Z => n337);
   U373 : CLKBUF_X1 port map( A => n393_port, Z => n338);
   U374 : CLKBUF_X1 port map( A => n393_port, Z => n339);
   U375 : CLKBUF_X1 port map( A => n393_port, Z => n340);
   U376 : CLKBUF_X1 port map( A => n393_port, Z => n341);
   U377 : CLKBUF_X1 port map( A => n393_port, Z => n342);
   U378 : CLKBUF_X1 port map( A => n393_port, Z => n343);
   U379 : CLKBUF_X1 port map( A => n392_port, Z => n344);
   U380 : CLKBUF_X1 port map( A => n392_port, Z => n345);
   U381 : CLKBUF_X1 port map( A => n392_port, Z => n346);
   U382 : CLKBUF_X1 port map( A => n392_port, Z => n347);
   U383 : CLKBUF_X1 port map( A => n392_port, Z => n348);
   U384 : CLKBUF_X1 port map( A => n392_port, Z => n349);
   U385 : CLKBUF_X1 port map( A => n391_port, Z => n350);
   U386 : CLKBUF_X1 port map( A => n391_port, Z => n351);
   U387 : CLKBUF_X1 port map( A => n391_port, Z => n352);
   U388 : CLKBUF_X1 port map( A => n391_port, Z => n353);
   U389 : CLKBUF_X1 port map( A => n391_port, Z => n354);
   U390 : CLKBUF_X1 port map( A => n391_port, Z => n355);
   U391 : CLKBUF_X1 port map( A => n390_port, Z => n356);
   U392 : CLKBUF_X1 port map( A => n390_port, Z => n357);
   U393 : CLKBUF_X1 port map( A => n390_port, Z => n358);
   U394 : CLKBUF_X1 port map( A => n390_port, Z => n359);
   U395 : CLKBUF_X1 port map( A => n390_port, Z => n360);
   U396 : CLKBUF_X1 port map( A => n390_port, Z => n361);
   U397 : CLKBUF_X1 port map( A => n389_port, Z => n362);
   U398 : CLKBUF_X1 port map( A => n389_port, Z => n363);
   U399 : CLKBUF_X1 port map( A => n389_port, Z => n364);
   U400 : CLKBUF_X1 port map( A => n389_port, Z => n365);
   U401 : CLKBUF_X1 port map( A => n389_port, Z => n366);
   U402 : CLKBUF_X1 port map( A => n389_port, Z => n367);
   U403 : CLKBUF_X1 port map( A => n388_port, Z => n368);
   U404 : CLKBUF_X1 port map( A => n388_port, Z => n369);
   U405 : CLKBUF_X1 port map( A => n388_port, Z => n370);
   U406 : CLKBUF_X1 port map( A => n388_port, Z => n371);
   U407 : CLKBUF_X1 port map( A => n388_port, Z => n372);
   U408 : CLKBUF_X1 port map( A => n388_port, Z => n373);
   U409 : CLKBUF_X1 port map( A => n387_port, Z => n374);
   U410 : CLKBUF_X1 port map( A => n387_port, Z => n375);
   U411 : CLKBUF_X1 port map( A => n387_port, Z => n376);
   U412 : CLKBUF_X1 port map( A => n387_port, Z => n377);
   U413 : CLKBUF_X1 port map( A => n387_port, Z => n378);
   U414 : CLKBUF_X1 port map( A => n387_port, Z => n379);
   U415 : CLKBUF_X1 port map( A => n386_port, Z => n380);
   U416 : CLKBUF_X1 port map( A => n386_port, Z => n381);
   U417 : CLKBUF_X1 port map( A => n386_port, Z => n382);
   U418 : CLKBUF_X1 port map( A => n386_port, Z => n383);
   U419 : CLKBUF_X1 port map( A => n386_port, Z => n384);
   U420 : CLKBUF_X1 port map( A => n386_port, Z => n385_port);
   U421 : NOR2_X1 port map( A1 => n1092, A2 => ADD_RD1(1), ZN => n403_port);
   U422 : AND2_X1 port map( A1 => n403_port, A2 => ADD_RD1(0), ZN => n1071);
   U423 : NOR2_X1 port map( A1 => n1092, A2 => n1093, ZN => n404_port);
   U424 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n404_port, ZN => n1070);
   U425 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n80, B1 => 
                           REGISTERS_23_0_port, B2 => n67, ZN => n410_port);
   U426 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n405_port
                           );
   U427 : AND2_X1 port map( A1 => n405_port, A2 => ADD_RD1(0), ZN => n1073);
   U428 : NOR2_X1 port map( A1 => n1093, A2 => ADD_RD1(2), ZN => n406_port);
   U429 : AND2_X1 port map( A1 => n406_port, A2 => ADD_RD1(0), ZN => n1072);
   U430 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n106_port, B1 => 
                           REGISTERS_19_0_port, B2 => n93, ZN => n409_port);
   U431 : AND2_X1 port map( A1 => n403_port, A2 => n1094, ZN => n1075);
   U432 : AND2_X1 port map( A1 => n404_port, A2 => n1094, ZN => n1074);
   U433 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n132, B1 => 
                           REGISTERS_22_0_port, B2 => n119_port, ZN => 
                           n408_port);
   U434 : AND2_X1 port map( A1 => n405_port, A2 => n1094, ZN => n1077);
   U435 : AND2_X1 port map( A1 => n406_port, A2 => n1094, ZN => n1076);
   U436 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n158, B1 => 
                           REGISTERS_18_0_port, B2 => n145, ZN => n407_port);
   U437 : AND4_X1 port map( A1 => n410_port, A2 => n409_port, A3 => n408_port, 
                           A4 => n407_port, ZN => n427_port);
   U438 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n80, B1 => 
                           REGISTERS_31_0_port, B2 => n67, ZN => n414_port);
   U439 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n106_port, B1 => 
                           REGISTERS_27_0_port, B2 => n93, ZN => n413_port);
   U440 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n132, B1 => 
                           REGISTERS_30_0_port, B2 => n119_port, ZN => 
                           n412_port);
   U441 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n158, B1 => 
                           REGISTERS_26_0_port, B2 => n145, ZN => n411_port);
   U442 : AND4_X1 port map( A1 => n414_port, A2 => n413_port, A3 => n412_port, 
                           A4 => n411_port, ZN => n426_port);
   U443 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n80, B1 => 
                           REGISTERS_7_0_port, B2 => n67, ZN => n418_port);
   U444 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n106_port, B1 => 
                           REGISTERS_3_0_port, B2 => n93, ZN => n417_port);
   U445 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n132, B1 => 
                           REGISTERS_6_0_port, B2 => n119_port, ZN => n416_port
                           );
   U446 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n158, B1 => 
                           REGISTERS_2_0_port, B2 => n145, ZN => n415_port);
   U447 : NAND4_X1 port map( A1 => n418_port, A2 => n417_port, A3 => n416_port,
                           A4 => n415_port, ZN => n424_port);
   U448 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n80, B1 => 
                           REGISTERS_15_0_port, B2 => n67, ZN => n422_port);
   U449 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n106_port, B1 => 
                           REGISTERS_11_0_port, B2 => n93, ZN => n421_port);
   U450 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n132, B1 => 
                           REGISTERS_14_0_port, B2 => n119_port, ZN => 
                           n420_port);
   U451 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n158, B1 => 
                           REGISTERS_10_0_port, B2 => n145, ZN => n419_port);
   U452 : NAND4_X1 port map( A1 => n422_port, A2 => n421_port, A3 => n420_port,
                           A4 => n419_port, ZN => n423_port);
   U453 : AOI22_X1 port map( A1 => n424_port, A2 => n1085, B1 => n423_port, B2 
                           => n1083, ZN => n425_port);
   U454 : OAI221_X1 port map( B1 => n1089, B2 => n427_port, C1 => n1087, C2 => 
                           n426_port, A => n425_port, ZN => N62);
   U455 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n80, B1 => 
                           REGISTERS_23_1_port, B2 => n67, ZN => n431_port);
   U456 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n106_port, B1 => 
                           REGISTERS_19_1_port, B2 => n93, ZN => n430_port);
   U457 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n132, B1 => 
                           REGISTERS_22_1_port, B2 => n119_port, ZN => 
                           n429_port);
   U458 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n158, B1 => 
                           REGISTERS_18_1_port, B2 => n145, ZN => n428_port);
   U459 : AND4_X1 port map( A1 => n431_port, A2 => n430_port, A3 => n429_port, 
                           A4 => n428_port, ZN => n448_port);
   U460 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n80, B1 => 
                           REGISTERS_31_1_port, B2 => n67, ZN => n435_port);
   U461 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n106_port, B1 => 
                           REGISTERS_27_1_port, B2 => n93, ZN => n434_port);
   U462 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n132, B1 => 
                           REGISTERS_30_1_port, B2 => n119_port, ZN => 
                           n433_port);
   U463 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n158, B1 => 
                           REGISTERS_26_1_port, B2 => n145, ZN => n432_port);
   U464 : AND4_X1 port map( A1 => n435_port, A2 => n434_port, A3 => n433_port, 
                           A4 => n432_port, ZN => n447_port);
   U465 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n80, B1 => 
                           REGISTERS_7_1_port, B2 => n67, ZN => n439_port);
   U466 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n106_port, B1 => 
                           REGISTERS_3_1_port, B2 => n93, ZN => n438_port);
   U467 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n132, B1 => 
                           REGISTERS_6_1_port, B2 => n119_port, ZN => n437_port
                           );
   U468 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n158, B1 => 
                           REGISTERS_2_1_port, B2 => n145, ZN => n436_port);
   U469 : NAND4_X1 port map( A1 => n439_port, A2 => n438_port, A3 => n437_port,
                           A4 => n436_port, ZN => n445_port);
   U470 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n80, B1 => 
                           REGISTERS_15_1_port, B2 => n67, ZN => n443_port);
   U471 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n106_port, B1 => 
                           REGISTERS_11_1_port, B2 => n93, ZN => n442_port);
   U472 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n132, B1 => 
                           REGISTERS_14_1_port, B2 => n119_port, ZN => 
                           n441_port);
   U473 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n158, B1 => 
                           REGISTERS_10_1_port, B2 => n145, ZN => n440_port);
   U474 : NAND4_X1 port map( A1 => n443_port, A2 => n442_port, A3 => n441_port,
                           A4 => n440_port, ZN => n444_port);
   U475 : AOI22_X1 port map( A1 => n445_port, A2 => n1085, B1 => n444_port, B2 
                           => n1083, ZN => n446_port);
   U476 : OAI221_X1 port map( B1 => n1089, B2 => n448_port, C1 => n1087, C2 => 
                           n447_port, A => n446_port, ZN => N61);
   U477 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n80, B1 => 
                           REGISTERS_23_2_port, B2 => n67, ZN => n452);
   U478 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n106_port, B1 => 
                           REGISTERS_19_2_port, B2 => n93, ZN => n451);
   U479 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n132, B1 => 
                           REGISTERS_22_2_port, B2 => n119_port, ZN => n450);
   U480 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n158, B1 => 
                           REGISTERS_18_2_port, B2 => n145, ZN => n449);
   U481 : AND4_X1 port map( A1 => n452, A2 => n451, A3 => n450, A4 => n449, ZN 
                           => n469);
   U482 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n80, B1 => 
                           REGISTERS_31_2_port, B2 => n67, ZN => n456);
   U483 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n106_port, B1 => 
                           REGISTERS_27_2_port, B2 => n93, ZN => n455);
   U484 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n132, B1 => 
                           REGISTERS_30_2_port, B2 => n119_port, ZN => n454);
   U485 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n158, B1 => 
                           REGISTERS_26_2_port, B2 => n145, ZN => n453);
   U486 : AND4_X1 port map( A1 => n456, A2 => n455, A3 => n454, A4 => n453, ZN 
                           => n468);
   U487 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n80, B1 => 
                           REGISTERS_7_2_port, B2 => n67, ZN => n460);
   U488 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n106_port, B1 => 
                           REGISTERS_3_2_port, B2 => n93, ZN => n459);
   U489 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n132, B1 => 
                           REGISTERS_6_2_port, B2 => n119_port, ZN => n458);
   U490 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n158, B1 => 
                           REGISTERS_2_2_port, B2 => n145, ZN => n457);
   U491 : NAND4_X1 port map( A1 => n460, A2 => n459, A3 => n458, A4 => n457, ZN
                           => n466);
   U492 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n80, B1 => 
                           REGISTERS_15_2_port, B2 => n67, ZN => n464);
   U493 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n106_port, B1 => 
                           REGISTERS_11_2_port, B2 => n93, ZN => n463);
   U494 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n132, B1 => 
                           REGISTERS_14_2_port, B2 => n119_port, ZN => n462);
   U495 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n158, B1 => 
                           REGISTERS_10_2_port, B2 => n145, ZN => n461);
   U496 : NAND4_X1 port map( A1 => n464, A2 => n463, A3 => n462, A4 => n461, ZN
                           => n465);
   U497 : AOI22_X1 port map( A1 => n466, A2 => n1085, B1 => n465, B2 => n1083, 
                           ZN => n467);
   U498 : OAI221_X1 port map( B1 => n1089, B2 => n469, C1 => n1087, C2 => n468,
                           A => n467, ZN => N60);
   U499 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n81, B1 => 
                           REGISTERS_23_3_port, B2 => n68, ZN => n473);
   U500 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n107_port, B1 => 
                           REGISTERS_19_3_port, B2 => n94, ZN => n472);
   U501 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n133, B1 => 
                           REGISTERS_22_3_port, B2 => n120_port, ZN => n471);
   U502 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n159, B1 => 
                           REGISTERS_18_3_port, B2 => n146, ZN => n470);
   U503 : AND4_X1 port map( A1 => n473, A2 => n472, A3 => n471, A4 => n470, ZN 
                           => n490);
   U504 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n81, B1 => 
                           REGISTERS_31_3_port, B2 => n68, ZN => n477);
   U505 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n107_port, B1 => 
                           REGISTERS_27_3_port, B2 => n94, ZN => n476);
   U506 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n133, B1 => 
                           REGISTERS_30_3_port, B2 => n120_port, ZN => n475);
   U507 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n159, B1 => 
                           REGISTERS_26_3_port, B2 => n146, ZN => n474);
   U508 : AND4_X1 port map( A1 => n477, A2 => n476, A3 => n475, A4 => n474, ZN 
                           => n489);
   U509 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n81, B1 => 
                           REGISTERS_7_3_port, B2 => n68, ZN => n481);
   U510 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n107_port, B1 => 
                           REGISTERS_3_3_port, B2 => n94, ZN => n480);
   U511 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n133, B1 => 
                           REGISTERS_6_3_port, B2 => n120_port, ZN => n479);
   U512 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n159, B1 => 
                           REGISTERS_2_3_port, B2 => n146, ZN => n478);
   U513 : NAND4_X1 port map( A1 => n481, A2 => n480, A3 => n479, A4 => n478, ZN
                           => n487);
   U514 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n81, B1 => 
                           REGISTERS_15_3_port, B2 => n68, ZN => n485);
   U515 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n107_port, B1 => 
                           REGISTERS_11_3_port, B2 => n94, ZN => n484);
   U516 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n133, B1 => 
                           REGISTERS_14_3_port, B2 => n120_port, ZN => n483);
   U517 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n159, B1 => 
                           REGISTERS_10_3_port, B2 => n146, ZN => n482);
   U518 : NAND4_X1 port map( A1 => n485, A2 => n484, A3 => n483, A4 => n482, ZN
                           => n486);
   U519 : AOI22_X1 port map( A1 => n487, A2 => n1085, B1 => n486, B2 => n1083, 
                           ZN => n488);
   U520 : OAI221_X1 port map( B1 => n1089, B2 => n490, C1 => n1087, C2 => n489,
                           A => n488, ZN => N59);
   U521 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n81, B1 => 
                           REGISTERS_23_4_port, B2 => n68, ZN => n494);
   U522 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n107_port, B1 => 
                           REGISTERS_19_4_port, B2 => n94, ZN => n493);
   U523 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n133, B1 => 
                           REGISTERS_22_4_port, B2 => n120_port, ZN => n492);
   U524 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n159, B1 => 
                           REGISTERS_18_4_port, B2 => n146, ZN => n491);
   U525 : AND4_X1 port map( A1 => n494, A2 => n493, A3 => n492, A4 => n491, ZN 
                           => n511);
   U526 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n81, B1 => 
                           REGISTERS_31_4_port, B2 => n68, ZN => n498);
   U527 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n107_port, B1 => 
                           REGISTERS_27_4_port, B2 => n94, ZN => n497);
   U528 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n133, B1 => 
                           REGISTERS_30_4_port, B2 => n120_port, ZN => n496);
   U529 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n159, B1 => 
                           REGISTERS_26_4_port, B2 => n146, ZN => n495);
   U530 : AND4_X1 port map( A1 => n498, A2 => n497, A3 => n496, A4 => n495, ZN 
                           => n510);
   U531 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n81, B1 => 
                           REGISTERS_7_4_port, B2 => n68, ZN => n502);
   U532 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n107_port, B1 => 
                           REGISTERS_3_4_port, B2 => n94, ZN => n501);
   U533 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n133, B1 => 
                           REGISTERS_6_4_port, B2 => n120_port, ZN => n500);
   U534 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n159, B1 => 
                           REGISTERS_2_4_port, B2 => n146, ZN => n499);
   U535 : NAND4_X1 port map( A1 => n502, A2 => n501, A3 => n500, A4 => n499, ZN
                           => n508);
   U536 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n81, B1 => 
                           REGISTERS_15_4_port, B2 => n68, ZN => n506);
   U537 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n107_port, B1 => 
                           REGISTERS_11_4_port, B2 => n94, ZN => n505);
   U538 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n133, B1 => 
                           REGISTERS_14_4_port, B2 => n120_port, ZN => n504);
   U539 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n159, B1 => 
                           REGISTERS_10_4_port, B2 => n146, ZN => n503);
   U540 : NAND4_X1 port map( A1 => n506, A2 => n505, A3 => n504, A4 => n503, ZN
                           => n507);
   U541 : AOI22_X1 port map( A1 => n508, A2 => n1085, B1 => n507, B2 => n1083, 
                           ZN => n509);
   U542 : OAI221_X1 port map( B1 => n1089, B2 => n511, C1 => n1087, C2 => n510,
                           A => n509, ZN => N58);
   U543 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n81, B1 => 
                           REGISTERS_23_5_port, B2 => n68, ZN => n515);
   U544 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n107_port, B1 => 
                           REGISTERS_19_5_port, B2 => n94, ZN => n514);
   U545 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n133, B1 => 
                           REGISTERS_22_5_port, B2 => n120_port, ZN => n513);
   U546 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n159, B1 => 
                           REGISTERS_18_5_port, B2 => n146, ZN => n512);
   U547 : AND4_X1 port map( A1 => n515, A2 => n514, A3 => n513, A4 => n512, ZN 
                           => n532);
   U548 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n81, B1 => 
                           REGISTERS_31_5_port, B2 => n68, ZN => n519);
   U549 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n107_port, B1 => 
                           REGISTERS_27_5_port, B2 => n94, ZN => n518);
   U550 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n133, B1 => 
                           REGISTERS_30_5_port, B2 => n120_port, ZN => n517);
   U551 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n159, B1 => 
                           REGISTERS_26_5_port, B2 => n146, ZN => n516);
   U552 : AND4_X1 port map( A1 => n519, A2 => n518, A3 => n517, A4 => n516, ZN 
                           => n531);
   U553 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n81, B1 => 
                           REGISTERS_7_5_port, B2 => n68, ZN => n523);
   U554 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n107_port, B1 => 
                           REGISTERS_3_5_port, B2 => n94, ZN => n522);
   U555 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n133, B1 => 
                           REGISTERS_6_5_port, B2 => n120_port, ZN => n521);
   U556 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n159, B1 => 
                           REGISTERS_2_5_port, B2 => n146, ZN => n520);
   U557 : NAND4_X1 port map( A1 => n523, A2 => n522, A3 => n521, A4 => n520, ZN
                           => n529);
   U558 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n81, B1 => 
                           REGISTERS_15_5_port, B2 => n68, ZN => n527);
   U559 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n107_port, B1 => 
                           REGISTERS_11_5_port, B2 => n94, ZN => n526);
   U560 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n133, B1 => 
                           REGISTERS_14_5_port, B2 => n120_port, ZN => n525);
   U561 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n159, B1 => 
                           REGISTERS_10_5_port, B2 => n146, ZN => n524);
   U562 : NAND4_X1 port map( A1 => n527, A2 => n526, A3 => n525, A4 => n524, ZN
                           => n528);
   U563 : AOI22_X1 port map( A1 => n529, A2 => n1085, B1 => n528, B2 => n1083, 
                           ZN => n530);
   U564 : OAI221_X1 port map( B1 => n1089, B2 => n532, C1 => n1087, C2 => n531,
                           A => n530, ZN => N57);
   U565 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n82, B1 => 
                           REGISTERS_23_6_port, B2 => n69, ZN => n536);
   U566 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n108_port, B1 => 
                           REGISTERS_19_6_port, B2 => n95, ZN => n535);
   U567 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n134, B1 => 
                           REGISTERS_22_6_port, B2 => n121_port, ZN => n534);
   U568 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n160, B1 => 
                           REGISTERS_18_6_port, B2 => n147, ZN => n533);
   U569 : AND4_X1 port map( A1 => n536, A2 => n535, A3 => n534, A4 => n533, ZN 
                           => n553);
   U570 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n82, B1 => 
                           REGISTERS_31_6_port, B2 => n69, ZN => n540);
   U571 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n108_port, B1 => 
                           REGISTERS_27_6_port, B2 => n95, ZN => n539);
   U572 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n134, B1 => 
                           REGISTERS_30_6_port, B2 => n121_port, ZN => n538);
   U573 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n160, B1 => 
                           REGISTERS_26_6_port, B2 => n147, ZN => n537);
   U574 : AND4_X1 port map( A1 => n540, A2 => n539, A3 => n538, A4 => n537, ZN 
                           => n552);
   U575 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n82, B1 => 
                           REGISTERS_7_6_port, B2 => n69, ZN => n544);
   U576 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n108_port, B1 => 
                           REGISTERS_3_6_port, B2 => n95, ZN => n543);
   U577 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n134, B1 => 
                           REGISTERS_6_6_port, B2 => n121_port, ZN => n542);
   U578 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n160, B1 => 
                           REGISTERS_2_6_port, B2 => n147, ZN => n541);
   U579 : NAND4_X1 port map( A1 => n544, A2 => n543, A3 => n542, A4 => n541, ZN
                           => n550);
   U580 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n82, B1 => 
                           REGISTERS_15_6_port, B2 => n69, ZN => n548);
   U581 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n108_port, B1 => 
                           REGISTERS_11_6_port, B2 => n95, ZN => n547);
   U582 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n134, B1 => 
                           REGISTERS_14_6_port, B2 => n121_port, ZN => n546);
   U583 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n160, B1 => 
                           REGISTERS_10_6_port, B2 => n147, ZN => n545);
   U584 : NAND4_X1 port map( A1 => n548, A2 => n547, A3 => n546, A4 => n545, ZN
                           => n549);
   U585 : AOI22_X1 port map( A1 => n550, A2 => n1085, B1 => n549, B2 => n1083, 
                           ZN => n551);
   U586 : OAI221_X1 port map( B1 => n1089, B2 => n553, C1 => n1087, C2 => n552,
                           A => n551, ZN => N56);
   U587 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n82, B1 => 
                           REGISTERS_23_7_port, B2 => n69, ZN => n557);
   U588 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n108_port, B1 => 
                           REGISTERS_19_7_port, B2 => n95, ZN => n556);
   U589 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n134, B1 => 
                           REGISTERS_22_7_port, B2 => n121_port, ZN => n555);
   U590 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n160, B1 => 
                           REGISTERS_18_7_port, B2 => n147, ZN => n554);
   U591 : AND4_X1 port map( A1 => n557, A2 => n556, A3 => n555, A4 => n554, ZN 
                           => n574);
   U592 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n82, B1 => 
                           REGISTERS_31_7_port, B2 => n69, ZN => n561);
   U593 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n108_port, B1 => 
                           REGISTERS_27_7_port, B2 => n95, ZN => n560);
   U594 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n134, B1 => 
                           REGISTERS_30_7_port, B2 => n121_port, ZN => n559);
   U595 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n160, B1 => 
                           REGISTERS_26_7_port, B2 => n147, ZN => n558);
   U596 : AND4_X1 port map( A1 => n561, A2 => n560, A3 => n559, A4 => n558, ZN 
                           => n573);
   U597 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n82, B1 => 
                           REGISTERS_7_7_port, B2 => n69, ZN => n565);
   U598 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n108_port, B1 => 
                           REGISTERS_3_7_port, B2 => n95, ZN => n564);
   U599 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n134, B1 => 
                           REGISTERS_6_7_port, B2 => n121_port, ZN => n563);
   U600 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n160, B1 => 
                           REGISTERS_2_7_port, B2 => n147, ZN => n562);
   U601 : NAND4_X1 port map( A1 => n565, A2 => n564, A3 => n563, A4 => n562, ZN
                           => n571);
   U602 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n82, B1 => 
                           REGISTERS_15_7_port, B2 => n69, ZN => n569);
   U603 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n108_port, B1 => 
                           REGISTERS_11_7_port, B2 => n95, ZN => n568);
   U604 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n134, B1 => 
                           REGISTERS_14_7_port, B2 => n121_port, ZN => n567);
   U605 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n160, B1 => 
                           REGISTERS_10_7_port, B2 => n147, ZN => n566);
   U606 : NAND4_X1 port map( A1 => n569, A2 => n568, A3 => n567, A4 => n566, ZN
                           => n570);
   U607 : AOI22_X1 port map( A1 => n571, A2 => n1085, B1 => n570, B2 => n1083, 
                           ZN => n572);
   U608 : OAI221_X1 port map( B1 => n1089, B2 => n574, C1 => n1087, C2 => n573,
                           A => n572, ZN => N55);
   U609 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n82, B1 => 
                           REGISTERS_23_8_port, B2 => n69, ZN => n578);
   U610 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n108_port, B1 => 
                           REGISTERS_19_8_port, B2 => n95, ZN => n577);
   U611 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n134, B1 => 
                           REGISTERS_22_8_port, B2 => n121_port, ZN => n576);
   U612 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n160, B1 => 
                           REGISTERS_18_8_port, B2 => n147, ZN => n575);
   U613 : AND4_X1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, ZN 
                           => n595);
   U614 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n82, B1 => 
                           REGISTERS_31_8_port, B2 => n69, ZN => n582);
   U615 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n108_port, B1 => 
                           REGISTERS_27_8_port, B2 => n95, ZN => n581);
   U616 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n134, B1 => 
                           REGISTERS_30_8_port, B2 => n121_port, ZN => n580);
   U617 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n160, B1 => 
                           REGISTERS_26_8_port, B2 => n147, ZN => n579);
   U618 : AND4_X1 port map( A1 => n582, A2 => n581, A3 => n580, A4 => n579, ZN 
                           => n594);
   U619 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n82, B1 => 
                           REGISTERS_7_8_port, B2 => n69, ZN => n586);
   U620 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n108_port, B1 => 
                           REGISTERS_3_8_port, B2 => n95, ZN => n585);
   U621 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n134, B1 => 
                           REGISTERS_6_8_port, B2 => n121_port, ZN => n584);
   U622 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n160, B1 => 
                           REGISTERS_2_8_port, B2 => n147, ZN => n583);
   U623 : NAND4_X1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, ZN
                           => n592);
   U624 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n82, B1 => 
                           REGISTERS_15_8_port, B2 => n69, ZN => n590);
   U625 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n108_port, B1 => 
                           REGISTERS_11_8_port, B2 => n95, ZN => n589);
   U626 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n134, B1 => 
                           REGISTERS_14_8_port, B2 => n121_port, ZN => n588);
   U627 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n160, B1 => 
                           REGISTERS_10_8_port, B2 => n147, ZN => n587);
   U628 : NAND4_X1 port map( A1 => n590, A2 => n589, A3 => n588, A4 => n587, ZN
                           => n591);
   U629 : AOI22_X1 port map( A1 => n592, A2 => n1085, B1 => n591, B2 => n1083, 
                           ZN => n593);
   U630 : OAI221_X1 port map( B1 => n1089, B2 => n595, C1 => n1087, C2 => n594,
                           A => n593, ZN => N54);
   U631 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n83, B1 => 
                           REGISTERS_23_9_port, B2 => n70, ZN => n599);
   U632 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n109_port, B1 => 
                           REGISTERS_19_9_port, B2 => n96_port, ZN => n598);
   U633 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n135, B1 => 
                           REGISTERS_22_9_port, B2 => n122_port, ZN => n597);
   U634 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n161, B1 => 
                           REGISTERS_18_9_port, B2 => n148, ZN => n596);
   U635 : AND4_X1 port map( A1 => n599, A2 => n598, A3 => n597, A4 => n596, ZN 
                           => n616);
   U636 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n83, B1 => 
                           REGISTERS_31_9_port, B2 => n70, ZN => n603);
   U637 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n109_port, B1 => 
                           REGISTERS_27_9_port, B2 => n96_port, ZN => n602);
   U638 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n135, B1 => 
                           REGISTERS_30_9_port, B2 => n122_port, ZN => n601);
   U639 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n161, B1 => 
                           REGISTERS_26_9_port, B2 => n148, ZN => n600);
   U640 : AND4_X1 port map( A1 => n603, A2 => n602, A3 => n601, A4 => n600, ZN 
                           => n615);
   U641 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n83, B1 => 
                           REGISTERS_7_9_port, B2 => n70, ZN => n607);
   U642 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n109_port, B1 => 
                           REGISTERS_3_9_port, B2 => n96_port, ZN => n606);
   U643 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n135, B1 => 
                           REGISTERS_6_9_port, B2 => n122_port, ZN => n605);
   U644 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n161, B1 => 
                           REGISTERS_2_9_port, B2 => n148, ZN => n604);
   U645 : NAND4_X1 port map( A1 => n607, A2 => n606, A3 => n605, A4 => n604, ZN
                           => n613);
   U646 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n83, B1 => 
                           REGISTERS_15_9_port, B2 => n70, ZN => n611);
   U647 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n109_port, B1 => 
                           REGISTERS_11_9_port, B2 => n96_port, ZN => n610);
   U648 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n135, B1 => 
                           REGISTERS_14_9_port, B2 => n122_port, ZN => n609);
   U649 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n161, B1 => 
                           REGISTERS_10_9_port, B2 => n148, ZN => n608);
   U650 : NAND4_X1 port map( A1 => n611, A2 => n610, A3 => n609, A4 => n608, ZN
                           => n612);
   U651 : AOI22_X1 port map( A1 => n613, A2 => n1085, B1 => n612, B2 => n1083, 
                           ZN => n614);
   U652 : OAI221_X1 port map( B1 => n1089, B2 => n616, C1 => n1087, C2 => n615,
                           A => n614, ZN => N53);
   U653 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n83, B1 => 
                           REGISTERS_23_10_port, B2 => n70, ZN => n620);
   U654 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n109_port, B1 =>
                           REGISTERS_19_10_port, B2 => n96_port, ZN => n619);
   U655 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n135, B1 => 
                           REGISTERS_22_10_port, B2 => n122_port, ZN => n618);
   U656 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n161, B1 => 
                           REGISTERS_18_10_port, B2 => n148, ZN => n617);
   U657 : AND4_X1 port map( A1 => n620, A2 => n619, A3 => n618, A4 => n617, ZN 
                           => n637);
   U658 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n83, B1 => 
                           REGISTERS_31_10_port, B2 => n70, ZN => n624);
   U659 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n109_port, B1 =>
                           REGISTERS_27_10_port, B2 => n96_port, ZN => n623);
   U660 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n135, B1 => 
                           REGISTERS_30_10_port, B2 => n122_port, ZN => n622);
   U661 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n161, B1 => 
                           REGISTERS_26_10_port, B2 => n148, ZN => n621);
   U662 : AND4_X1 port map( A1 => n624, A2 => n623, A3 => n622, A4 => n621, ZN 
                           => n636);
   U663 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n83, B1 => 
                           REGISTERS_7_10_port, B2 => n70, ZN => n628);
   U664 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n109_port, B1 => 
                           REGISTERS_3_10_port, B2 => n96_port, ZN => n627);
   U665 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n135, B1 => 
                           REGISTERS_6_10_port, B2 => n122_port, ZN => n626);
   U666 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n161, B1 => 
                           REGISTERS_2_10_port, B2 => n148, ZN => n625);
   U667 : NAND4_X1 port map( A1 => n628, A2 => n627, A3 => n626, A4 => n625, ZN
                           => n634);
   U668 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n83, B1 => 
                           REGISTERS_15_10_port, B2 => n70, ZN => n632);
   U669 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n109_port, B1 => 
                           REGISTERS_11_10_port, B2 => n96_port, ZN => n631);
   U670 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n135, B1 => 
                           REGISTERS_14_10_port, B2 => n122_port, ZN => n630);
   U671 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n161, B1 => 
                           REGISTERS_10_10_port, B2 => n148, ZN => n629);
   U672 : NAND4_X1 port map( A1 => n632, A2 => n631, A3 => n630, A4 => n629, ZN
                           => n633);
   U673 : AOI22_X1 port map( A1 => n634, A2 => n1085, B1 => n633, B2 => n1083, 
                           ZN => n635);
   U674 : OAI221_X1 port map( B1 => n1089, B2 => n637, C1 => n1087, C2 => n636,
                           A => n635, ZN => N52);
   U675 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n83, B1 => 
                           REGISTERS_23_11_port, B2 => n70, ZN => n641);
   U676 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n109_port, B1 =>
                           REGISTERS_19_11_port, B2 => n96_port, ZN => n640);
   U677 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n135, B1 => 
                           REGISTERS_22_11_port, B2 => n122_port, ZN => n639);
   U678 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n161, B1 => 
                           REGISTERS_18_11_port, B2 => n148, ZN => n638);
   U679 : AND4_X1 port map( A1 => n641, A2 => n640, A3 => n639, A4 => n638, ZN 
                           => n658);
   U680 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n83, B1 => 
                           REGISTERS_31_11_port, B2 => n70, ZN => n645);
   U681 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n109_port, B1 =>
                           REGISTERS_27_11_port, B2 => n96_port, ZN => n644);
   U682 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n135, B1 => 
                           REGISTERS_30_11_port, B2 => n122_port, ZN => n643);
   U683 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n161, B1 => 
                           REGISTERS_26_11_port, B2 => n148, ZN => n642);
   U684 : AND4_X1 port map( A1 => n645, A2 => n644, A3 => n643, A4 => n642, ZN 
                           => n657);
   U685 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n83, B1 => 
                           REGISTERS_7_11_port, B2 => n70, ZN => n649);
   U686 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n109_port, B1 => 
                           REGISTERS_3_11_port, B2 => n96_port, ZN => n648);
   U687 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n135, B1 => 
                           REGISTERS_6_11_port, B2 => n122_port, ZN => n647);
   U688 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n161, B1 => 
                           REGISTERS_2_11_port, B2 => n148, ZN => n646);
   U689 : NAND4_X1 port map( A1 => n649, A2 => n648, A3 => n647, A4 => n646, ZN
                           => n655);
   U690 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n83, B1 => 
                           REGISTERS_15_11_port, B2 => n70, ZN => n653);
   U691 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n109_port, B1 => 
                           REGISTERS_11_11_port, B2 => n96_port, ZN => n652);
   U692 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n135, B1 => 
                           REGISTERS_14_11_port, B2 => n122_port, ZN => n651);
   U693 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n161, B1 => 
                           REGISTERS_10_11_port, B2 => n148, ZN => n650);
   U694 : NAND4_X1 port map( A1 => n653, A2 => n652, A3 => n651, A4 => n650, ZN
                           => n654);
   U695 : AOI22_X1 port map( A1 => n655, A2 => n1085, B1 => n654, B2 => n1083, 
                           ZN => n656);
   U696 : OAI221_X1 port map( B1 => n1089, B2 => n658, C1 => n1087, C2 => n657,
                           A => n656, ZN => N51);
   U697 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n84, B1 => 
                           REGISTERS_23_12_port, B2 => n71, ZN => n662);
   U698 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n110_port, B1 =>
                           REGISTERS_19_12_port, B2 => n97_port, ZN => n661);
   U699 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n136, B1 => 
                           REGISTERS_22_12_port, B2 => n123_port, ZN => n660);
   U700 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n162, B1 => 
                           REGISTERS_18_12_port, B2 => n149, ZN => n659);
   U701 : AND4_X1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, ZN 
                           => n679);
   U702 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n84, B1 => 
                           REGISTERS_31_12_port, B2 => n71, ZN => n666);
   U703 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n110_port, B1 =>
                           REGISTERS_27_12_port, B2 => n97_port, ZN => n665);
   U704 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n136, B1 => 
                           REGISTERS_30_12_port, B2 => n123_port, ZN => n664);
   U705 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n162, B1 => 
                           REGISTERS_26_12_port, B2 => n149, ZN => n663);
   U706 : AND4_X1 port map( A1 => n666, A2 => n665, A3 => n664, A4 => n663, ZN 
                           => n678);
   U707 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n84, B1 => 
                           REGISTERS_7_12_port, B2 => n71, ZN => n670);
   U708 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n110_port, B1 => 
                           REGISTERS_3_12_port, B2 => n97_port, ZN => n669);
   U709 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n136, B1 => 
                           REGISTERS_6_12_port, B2 => n123_port, ZN => n668);
   U710 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n162, B1 => 
                           REGISTERS_2_12_port, B2 => n149, ZN => n667);
   U711 : NAND4_X1 port map( A1 => n670, A2 => n669, A3 => n668, A4 => n667, ZN
                           => n676);
   U712 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n84, B1 => 
                           REGISTERS_15_12_port, B2 => n71, ZN => n674);
   U713 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n110_port, B1 => 
                           REGISTERS_11_12_port, B2 => n97_port, ZN => n673);
   U714 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n136, B1 => 
                           REGISTERS_14_12_port, B2 => n123_port, ZN => n672);
   U715 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n162, B1 => 
                           REGISTERS_10_12_port, B2 => n149, ZN => n671);
   U716 : NAND4_X1 port map( A1 => n674, A2 => n673, A3 => n672, A4 => n671, ZN
                           => n675);
   U717 : AOI22_X1 port map( A1 => n676, A2 => n1085, B1 => n675, B2 => n1083, 
                           ZN => n677);
   U718 : OAI221_X1 port map( B1 => n1089, B2 => n679, C1 => n1087, C2 => n678,
                           A => n677, ZN => N50);
   U719 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n84, B1 => 
                           REGISTERS_23_13_port, B2 => n71, ZN => n683);
   U720 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n110_port, B1 =>
                           REGISTERS_19_13_port, B2 => n97_port, ZN => n682);
   U721 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n136, B1 => 
                           REGISTERS_22_13_port, B2 => n123_port, ZN => n681);
   U722 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n162, B1 => 
                           REGISTERS_18_13_port, B2 => n149, ZN => n680);
   U723 : AND4_X1 port map( A1 => n683, A2 => n682, A3 => n681, A4 => n680, ZN 
                           => n700);
   U724 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n84, B1 => 
                           REGISTERS_31_13_port, B2 => n71, ZN => n687);
   U725 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n110_port, B1 =>
                           REGISTERS_27_13_port, B2 => n97_port, ZN => n686);
   U726 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n136, B1 => 
                           REGISTERS_30_13_port, B2 => n123_port, ZN => n685);
   U727 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n162, B1 => 
                           REGISTERS_26_13_port, B2 => n149, ZN => n684);
   U728 : AND4_X1 port map( A1 => n687, A2 => n686, A3 => n685, A4 => n684, ZN 
                           => n699);
   U729 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n84, B1 => 
                           REGISTERS_7_13_port, B2 => n71, ZN => n691);
   U730 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n110_port, B1 => 
                           REGISTERS_3_13_port, B2 => n97_port, ZN => n690);
   U731 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n136, B1 => 
                           REGISTERS_6_13_port, B2 => n123_port, ZN => n689);
   U732 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n162, B1 => 
                           REGISTERS_2_13_port, B2 => n149, ZN => n688);
   U733 : NAND4_X1 port map( A1 => n691, A2 => n690, A3 => n689, A4 => n688, ZN
                           => n697);
   U734 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n84, B1 => 
                           REGISTERS_15_13_port, B2 => n71, ZN => n695);
   U735 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n110_port, B1 => 
                           REGISTERS_11_13_port, B2 => n97_port, ZN => n694);
   U736 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n136, B1 => 
                           REGISTERS_14_13_port, B2 => n123_port, ZN => n693);
   U737 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n162, B1 => 
                           REGISTERS_10_13_port, B2 => n149, ZN => n692);
   U738 : NAND4_X1 port map( A1 => n695, A2 => n694, A3 => n693, A4 => n692, ZN
                           => n696);
   U739 : AOI22_X1 port map( A1 => n697, A2 => n1085, B1 => n696, B2 => n1083, 
                           ZN => n698);
   U740 : OAI221_X1 port map( B1 => n1089, B2 => n700, C1 => n1087, C2 => n699,
                           A => n698, ZN => N49);
   U741 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n84, B1 => 
                           REGISTERS_23_14_port, B2 => n71, ZN => n704);
   U742 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n110_port, B1 =>
                           REGISTERS_19_14_port, B2 => n97_port, ZN => n703);
   U743 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n136, B1 => 
                           REGISTERS_22_14_port, B2 => n123_port, ZN => n702);
   U744 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n162, B1 => 
                           REGISTERS_18_14_port, B2 => n149, ZN => n701);
   U745 : AND4_X1 port map( A1 => n704, A2 => n703, A3 => n702, A4 => n701, ZN 
                           => n721);
   U746 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n84, B1 => 
                           REGISTERS_31_14_port, B2 => n71, ZN => n708);
   U747 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n110_port, B1 =>
                           REGISTERS_27_14_port, B2 => n97_port, ZN => n707);
   U748 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n136, B1 => 
                           REGISTERS_30_14_port, B2 => n123_port, ZN => n706);
   U749 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n162, B1 => 
                           REGISTERS_26_14_port, B2 => n149, ZN => n705);
   U750 : AND4_X1 port map( A1 => n708, A2 => n707, A3 => n706, A4 => n705, ZN 
                           => n720);
   U751 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n84, B1 => 
                           REGISTERS_7_14_port, B2 => n71, ZN => n712);
   U752 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n110_port, B1 => 
                           REGISTERS_3_14_port, B2 => n97_port, ZN => n711);
   U753 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n136, B1 => 
                           REGISTERS_6_14_port, B2 => n123_port, ZN => n710);
   U754 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n162, B1 => 
                           REGISTERS_2_14_port, B2 => n149, ZN => n709);
   U755 : NAND4_X1 port map( A1 => n712, A2 => n711, A3 => n710, A4 => n709, ZN
                           => n718);
   U756 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n84, B1 => 
                           REGISTERS_15_14_port, B2 => n71, ZN => n716);
   U757 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n110_port, B1 => 
                           REGISTERS_11_14_port, B2 => n97_port, ZN => n715);
   U758 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n136, B1 => 
                           REGISTERS_14_14_port, B2 => n123_port, ZN => n714);
   U759 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n162, B1 => 
                           REGISTERS_10_14_port, B2 => n149, ZN => n713);
   U760 : NAND4_X1 port map( A1 => n716, A2 => n715, A3 => n714, A4 => n713, ZN
                           => n717);
   U761 : AOI22_X1 port map( A1 => n718, A2 => n1085, B1 => n717, B2 => n1083, 
                           ZN => n719);
   U762 : OAI221_X1 port map( B1 => n1089, B2 => n721, C1 => n1087, C2 => n720,
                           A => n719, ZN => N48);
   U763 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n85, B1 => 
                           REGISTERS_23_15_port, B2 => n72, ZN => n725);
   U764 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n111_port, B1 =>
                           REGISTERS_19_15_port, B2 => n98_port, ZN => n724);
   U765 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n137, B1 => 
                           REGISTERS_22_15_port, B2 => n124_port, ZN => n723);
   U766 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n163, B1 => 
                           REGISTERS_18_15_port, B2 => n150, ZN => n722);
   U767 : AND4_X1 port map( A1 => n725, A2 => n724, A3 => n723, A4 => n722, ZN 
                           => n742);
   U768 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n85, B1 => 
                           REGISTERS_31_15_port, B2 => n72, ZN => n729);
   U769 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n111_port, B1 =>
                           REGISTERS_27_15_port, B2 => n98_port, ZN => n728);
   U770 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n137, B1 => 
                           REGISTERS_30_15_port, B2 => n124_port, ZN => n727);
   U771 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n163, B1 => 
                           REGISTERS_26_15_port, B2 => n150, ZN => n726);
   U772 : AND4_X1 port map( A1 => n729, A2 => n728, A3 => n727, A4 => n726, ZN 
                           => n741);
   U773 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n85, B1 => 
                           REGISTERS_7_15_port, B2 => n72, ZN => n733);
   U774 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n111_port, B1 => 
                           REGISTERS_3_15_port, B2 => n98_port, ZN => n732);
   U775 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n137, B1 => 
                           REGISTERS_6_15_port, B2 => n124_port, ZN => n731);
   U776 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n163, B1 => 
                           REGISTERS_2_15_port, B2 => n150, ZN => n730);
   U777 : NAND4_X1 port map( A1 => n733, A2 => n732, A3 => n731, A4 => n730, ZN
                           => n739);
   U778 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n85, B1 => 
                           REGISTERS_15_15_port, B2 => n72, ZN => n737);
   U779 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n111_port, B1 => 
                           REGISTERS_11_15_port, B2 => n98_port, ZN => n736);
   U780 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n137, B1 => 
                           REGISTERS_14_15_port, B2 => n124_port, ZN => n735);
   U781 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n163, B1 => 
                           REGISTERS_10_15_port, B2 => n150, ZN => n734);
   U782 : NAND4_X1 port map( A1 => n737, A2 => n736, A3 => n735, A4 => n734, ZN
                           => n738);
   U783 : AOI22_X1 port map( A1 => n739, A2 => n1085, B1 => n738, B2 => n1083, 
                           ZN => n740);
   U784 : OAI221_X1 port map( B1 => n1089, B2 => n742, C1 => n1087, C2 => n741,
                           A => n740, ZN => N47);
   U785 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n85, B1 => 
                           REGISTERS_23_16_port, B2 => n72, ZN => n746);
   U786 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n111_port, B1 =>
                           REGISTERS_19_16_port, B2 => n98_port, ZN => n745);
   U787 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n137, B1 => 
                           REGISTERS_22_16_port, B2 => n124_port, ZN => n744);
   U788 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n163, B1 => 
                           REGISTERS_18_16_port, B2 => n150, ZN => n743);
   U789 : AND4_X1 port map( A1 => n746, A2 => n745, A3 => n744, A4 => n743, ZN 
                           => n763);
   U790 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n85, B1 => 
                           REGISTERS_31_16_port, B2 => n72, ZN => n750);
   U791 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n111_port, B1 =>
                           REGISTERS_27_16_port, B2 => n98_port, ZN => n749);
   U792 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n137, B1 => 
                           REGISTERS_30_16_port, B2 => n124_port, ZN => n748);
   U793 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n163, B1 => 
                           REGISTERS_26_16_port, B2 => n150, ZN => n747);
   U794 : AND4_X1 port map( A1 => n750, A2 => n749, A3 => n748, A4 => n747, ZN 
                           => n762);
   U795 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n85, B1 => 
                           REGISTERS_7_16_port, B2 => n72, ZN => n754);
   U796 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n111_port, B1 => 
                           REGISTERS_3_16_port, B2 => n98_port, ZN => n753);
   U797 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n137, B1 => 
                           REGISTERS_6_16_port, B2 => n124_port, ZN => n752);
   U798 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n163, B1 => 
                           REGISTERS_2_16_port, B2 => n150, ZN => n751);
   U799 : NAND4_X1 port map( A1 => n754, A2 => n753, A3 => n752, A4 => n751, ZN
                           => n760);
   U800 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n85, B1 => 
                           REGISTERS_15_16_port, B2 => n72, ZN => n758);
   U801 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n111_port, B1 => 
                           REGISTERS_11_16_port, B2 => n98_port, ZN => n757);
   U802 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n137, B1 => 
                           REGISTERS_14_16_port, B2 => n124_port, ZN => n756);
   U803 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n163, B1 => 
                           REGISTERS_10_16_port, B2 => n150, ZN => n755);
   U804 : NAND4_X1 port map( A1 => n758, A2 => n757, A3 => n756, A4 => n755, ZN
                           => n759);
   U805 : AOI22_X1 port map( A1 => n760, A2 => n1085, B1 => n759, B2 => n1083, 
                           ZN => n761);
   U806 : OAI221_X1 port map( B1 => n1089, B2 => n763, C1 => n1087, C2 => n762,
                           A => n761, ZN => N46);
   U807 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n85, B1 => 
                           REGISTERS_23_17_port, B2 => n72, ZN => n767);
   U808 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n111_port, B1 =>
                           REGISTERS_19_17_port, B2 => n98_port, ZN => n766);
   U809 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n137, B1 => 
                           REGISTERS_22_17_port, B2 => n124_port, ZN => n765);
   U810 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n163, B1 => 
                           REGISTERS_18_17_port, B2 => n150, ZN => n764);
   U811 : AND4_X1 port map( A1 => n767, A2 => n766, A3 => n765, A4 => n764, ZN 
                           => n784);
   U812 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n85, B1 => 
                           REGISTERS_31_17_port, B2 => n72, ZN => n771);
   U813 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n111_port, B1 =>
                           REGISTERS_27_17_port, B2 => n98_port, ZN => n770);
   U814 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n137, B1 => 
                           REGISTERS_30_17_port, B2 => n124_port, ZN => n769);
   U815 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n163, B1 => 
                           REGISTERS_26_17_port, B2 => n150, ZN => n768);
   U816 : AND4_X1 port map( A1 => n771, A2 => n770, A3 => n769, A4 => n768, ZN 
                           => n783);
   U817 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n85, B1 => 
                           REGISTERS_7_17_port, B2 => n72, ZN => n775);
   U818 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n111_port, B1 => 
                           REGISTERS_3_17_port, B2 => n98_port, ZN => n774);
   U819 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n137, B1 => 
                           REGISTERS_6_17_port, B2 => n124_port, ZN => n773);
   U820 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n163, B1 => 
                           REGISTERS_2_17_port, B2 => n150, ZN => n772);
   U821 : NAND4_X1 port map( A1 => n775, A2 => n774, A3 => n773, A4 => n772, ZN
                           => n781);
   U822 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n85, B1 => 
                           REGISTERS_15_17_port, B2 => n72, ZN => n779);
   U823 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n111_port, B1 => 
                           REGISTERS_11_17_port, B2 => n98_port, ZN => n778);
   U824 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n137, B1 => 
                           REGISTERS_14_17_port, B2 => n124_port, ZN => n777);
   U825 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n163, B1 => 
                           REGISTERS_10_17_port, B2 => n150, ZN => n776);
   U826 : NAND4_X1 port map( A1 => n779, A2 => n778, A3 => n777, A4 => n776, ZN
                           => n780);
   U827 : AOI22_X1 port map( A1 => n781, A2 => n1085, B1 => n780, B2 => n1083, 
                           ZN => n782);
   U828 : OAI221_X1 port map( B1 => n1089, B2 => n784, C1 => n1087, C2 => n783,
                           A => n782, ZN => N45);
   U829 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n86, B1 => 
                           REGISTERS_23_18_port, B2 => n73, ZN => n788);
   U830 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n112_port, B1 =>
                           REGISTERS_19_18_port, B2 => n99_port, ZN => n787);
   U831 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n138, B1 => 
                           REGISTERS_22_18_port, B2 => n125_port, ZN => n786);
   U832 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n164, B1 => 
                           REGISTERS_18_18_port, B2 => n151, ZN => n785);
   U833 : AND4_X1 port map( A1 => n788, A2 => n787, A3 => n786, A4 => n785, ZN 
                           => n805);
   U834 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n86, B1 => 
                           REGISTERS_31_18_port, B2 => n73, ZN => n792);
   U835 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n112_port, B1 =>
                           REGISTERS_27_18_port, B2 => n99_port, ZN => n791);
   U836 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n138, B1 => 
                           REGISTERS_30_18_port, B2 => n125_port, ZN => n790);
   U837 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n164, B1 => 
                           REGISTERS_26_18_port, B2 => n151, ZN => n789);
   U838 : AND4_X1 port map( A1 => n792, A2 => n791, A3 => n790, A4 => n789, ZN 
                           => n804);
   U839 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n86, B1 => 
                           REGISTERS_7_18_port, B2 => n73, ZN => n796);
   U840 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n112_port, B1 => 
                           REGISTERS_3_18_port, B2 => n99_port, ZN => n795);
   U841 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n138, B1 => 
                           REGISTERS_6_18_port, B2 => n125_port, ZN => n794);
   U842 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n164, B1 => 
                           REGISTERS_2_18_port, B2 => n151, ZN => n793);
   U843 : NAND4_X1 port map( A1 => n796, A2 => n795, A3 => n794, A4 => n793, ZN
                           => n802);
   U844 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n86, B1 => 
                           REGISTERS_15_18_port, B2 => n73, ZN => n800);
   U845 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n112_port, B1 => 
                           REGISTERS_11_18_port, B2 => n99_port, ZN => n799);
   U846 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n138, B1 => 
                           REGISTERS_14_18_port, B2 => n125_port, ZN => n798);
   U847 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n164, B1 => 
                           REGISTERS_10_18_port, B2 => n151, ZN => n797);
   U848 : NAND4_X1 port map( A1 => n800, A2 => n799, A3 => n798, A4 => n797, ZN
                           => n801);
   U849 : AOI22_X1 port map( A1 => n802, A2 => n1085, B1 => n801, B2 => n1083, 
                           ZN => n803);
   U850 : OAI221_X1 port map( B1 => n1089, B2 => n805, C1 => n1087, C2 => n804,
                           A => n803, ZN => N44);
   U851 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n86, B1 => 
                           REGISTERS_23_19_port, B2 => n73, ZN => n809);
   U852 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n112_port, B1 =>
                           REGISTERS_19_19_port, B2 => n99_port, ZN => n808);
   U853 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n138, B1 => 
                           REGISTERS_22_19_port, B2 => n125_port, ZN => n807);
   U854 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n164, B1 => 
                           REGISTERS_18_19_port, B2 => n151, ZN => n806);
   U855 : AND4_X1 port map( A1 => n809, A2 => n808, A3 => n807, A4 => n806, ZN 
                           => n826);
   U856 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n86, B1 => 
                           REGISTERS_31_19_port, B2 => n73, ZN => n813);
   U857 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n112_port, B1 =>
                           REGISTERS_27_19_port, B2 => n99_port, ZN => n812);
   U858 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n138, B1 => 
                           REGISTERS_30_19_port, B2 => n125_port, ZN => n811);
   U859 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n164, B1 => 
                           REGISTERS_26_19_port, B2 => n151, ZN => n810);
   U860 : AND4_X1 port map( A1 => n813, A2 => n812, A3 => n811, A4 => n810, ZN 
                           => n825);
   U861 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n86, B1 => 
                           REGISTERS_7_19_port, B2 => n73, ZN => n817);
   U862 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n112_port, B1 => 
                           REGISTERS_3_19_port, B2 => n99_port, ZN => n816);
   U863 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n138, B1 => 
                           REGISTERS_6_19_port, B2 => n125_port, ZN => n815);
   U864 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n164, B1 => 
                           REGISTERS_2_19_port, B2 => n151, ZN => n814);
   U865 : NAND4_X1 port map( A1 => n817, A2 => n816, A3 => n815, A4 => n814, ZN
                           => n823);
   U866 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n86, B1 => 
                           REGISTERS_15_19_port, B2 => n73, ZN => n821);
   U867 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n112_port, B1 => 
                           REGISTERS_11_19_port, B2 => n99_port, ZN => n820);
   U868 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n138, B1 => 
                           REGISTERS_14_19_port, B2 => n125_port, ZN => n819);
   U869 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n164, B1 => 
                           REGISTERS_10_19_port, B2 => n151, ZN => n818);
   U870 : NAND4_X1 port map( A1 => n821, A2 => n820, A3 => n819, A4 => n818, ZN
                           => n822);
   U871 : AOI22_X1 port map( A1 => n823, A2 => n1085, B1 => n822, B2 => n1083, 
                           ZN => n824);
   U872 : OAI221_X1 port map( B1 => n1089, B2 => n826, C1 => n1087, C2 => n825,
                           A => n824, ZN => N43);
   U873 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n86, B1 => 
                           REGISTERS_23_20_port, B2 => n73, ZN => n830);
   U874 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n112_port, B1 =>
                           REGISTERS_19_20_port, B2 => n99_port, ZN => n829);
   U875 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n138, B1 => 
                           REGISTERS_22_20_port, B2 => n125_port, ZN => n828);
   U876 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n164, B1 => 
                           REGISTERS_18_20_port, B2 => n151, ZN => n827);
   U877 : AND4_X1 port map( A1 => n830, A2 => n829, A3 => n828, A4 => n827, ZN 
                           => n847);
   U878 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n86, B1 => 
                           REGISTERS_31_20_port, B2 => n73, ZN => n834);
   U879 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n112_port, B1 =>
                           REGISTERS_27_20_port, B2 => n99_port, ZN => n833);
   U880 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n138, B1 => 
                           REGISTERS_30_20_port, B2 => n125_port, ZN => n832);
   U881 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n164, B1 => 
                           REGISTERS_26_20_port, B2 => n151, ZN => n831);
   U882 : AND4_X1 port map( A1 => n834, A2 => n833, A3 => n832, A4 => n831, ZN 
                           => n846);
   U883 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n86, B1 => 
                           REGISTERS_7_20_port, B2 => n73, ZN => n838);
   U884 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n112_port, B1 => 
                           REGISTERS_3_20_port, B2 => n99_port, ZN => n837);
   U885 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n138, B1 => 
                           REGISTERS_6_20_port, B2 => n125_port, ZN => n836);
   U886 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n164, B1 => 
                           REGISTERS_2_20_port, B2 => n151, ZN => n835);
   U887 : NAND4_X1 port map( A1 => n838, A2 => n837, A3 => n836, A4 => n835, ZN
                           => n844);
   U888 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n86, B1 => 
                           REGISTERS_15_20_port, B2 => n73, ZN => n842);
   U889 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n112_port, B1 => 
                           REGISTERS_11_20_port, B2 => n99_port, ZN => n841);
   U890 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n138, B1 => 
                           REGISTERS_14_20_port, B2 => n125_port, ZN => n840);
   U891 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n164, B1 => 
                           REGISTERS_10_20_port, B2 => n151, ZN => n839);
   U892 : NAND4_X1 port map( A1 => n842, A2 => n841, A3 => n840, A4 => n839, ZN
                           => n843);
   U893 : AOI22_X1 port map( A1 => n844, A2 => n1085, B1 => n843, B2 => n1083, 
                           ZN => n845);
   U894 : OAI221_X1 port map( B1 => n1089, B2 => n847, C1 => n1087, C2 => n846,
                           A => n845, ZN => N42);
   U895 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n87, B1 => 
                           REGISTERS_23_21_port, B2 => n74, ZN => n851);
   U896 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n113_port, B1 =>
                           REGISTERS_19_21_port, B2 => n100_port, ZN => n850);
   U897 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n139, B1 => 
                           REGISTERS_22_21_port, B2 => n126_port, ZN => n849);
   U898 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n165, B1 => 
                           REGISTERS_18_21_port, B2 => n152, ZN => n848);
   U899 : AND4_X1 port map( A1 => n851, A2 => n850, A3 => n849, A4 => n848, ZN 
                           => n868);
   U900 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n87, B1 => 
                           REGISTERS_31_21_port, B2 => n74, ZN => n855);
   U901 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n113_port, B1 =>
                           REGISTERS_27_21_port, B2 => n100_port, ZN => n854);
   U902 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n139, B1 => 
                           REGISTERS_30_21_port, B2 => n126_port, ZN => n853);
   U903 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n165, B1 => 
                           REGISTERS_26_21_port, B2 => n152, ZN => n852);
   U904 : AND4_X1 port map( A1 => n855, A2 => n854, A3 => n853, A4 => n852, ZN 
                           => n867);
   U905 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n87, B1 => 
                           REGISTERS_7_21_port, B2 => n74, ZN => n859);
   U906 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n113_port, B1 => 
                           REGISTERS_3_21_port, B2 => n100_port, ZN => n858);
   U907 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n139, B1 => 
                           REGISTERS_6_21_port, B2 => n126_port, ZN => n857);
   U908 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n165, B1 => 
                           REGISTERS_2_21_port, B2 => n152, ZN => n856);
   U909 : NAND4_X1 port map( A1 => n859, A2 => n858, A3 => n857, A4 => n856, ZN
                           => n865);
   U910 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n87, B1 => 
                           REGISTERS_15_21_port, B2 => n74, ZN => n863);
   U911 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n113_port, B1 => 
                           REGISTERS_11_21_port, B2 => n100_port, ZN => n862);
   U912 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n139, B1 => 
                           REGISTERS_14_21_port, B2 => n126_port, ZN => n861);
   U913 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n165, B1 => 
                           REGISTERS_10_21_port, B2 => n152, ZN => n860);
   U914 : NAND4_X1 port map( A1 => n863, A2 => n862, A3 => n861, A4 => n860, ZN
                           => n864);
   U915 : AOI22_X1 port map( A1 => n865, A2 => n1085, B1 => n864, B2 => n1083, 
                           ZN => n866);
   U916 : OAI221_X1 port map( B1 => n1089, B2 => n868, C1 => n1087, C2 => n867,
                           A => n866, ZN => N41);
   U917 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n87, B1 => 
                           REGISTERS_23_22_port, B2 => n74, ZN => n872);
   U918 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n113_port, B1 =>
                           REGISTERS_19_22_port, B2 => n100_port, ZN => n871);
   U919 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n139, B1 => 
                           REGISTERS_22_22_port, B2 => n126_port, ZN => n870);
   U920 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n165, B1 => 
                           REGISTERS_18_22_port, B2 => n152, ZN => n869);
   U921 : AND4_X1 port map( A1 => n872, A2 => n871, A3 => n870, A4 => n869, ZN 
                           => n889);
   U922 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n87, B1 => 
                           REGISTERS_31_22_port, B2 => n74, ZN => n876);
   U923 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n113_port, B1 =>
                           REGISTERS_27_22_port, B2 => n100_port, ZN => n875);
   U924 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n139, B1 => 
                           REGISTERS_30_22_port, B2 => n126_port, ZN => n874);
   U925 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n165, B1 => 
                           REGISTERS_26_22_port, B2 => n152, ZN => n873);
   U926 : AND4_X1 port map( A1 => n876, A2 => n875, A3 => n874, A4 => n873, ZN 
                           => n888);
   U927 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n87, B1 => 
                           REGISTERS_7_22_port, B2 => n74, ZN => n880);
   U928 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n113_port, B1 => 
                           REGISTERS_3_22_port, B2 => n100_port, ZN => n879);
   U929 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n139, B1 => 
                           REGISTERS_6_22_port, B2 => n126_port, ZN => n878);
   U930 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n165, B1 => 
                           REGISTERS_2_22_port, B2 => n152, ZN => n877);
   U931 : NAND4_X1 port map( A1 => n880, A2 => n879, A3 => n878, A4 => n877, ZN
                           => n886);
   U932 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n87, B1 => 
                           REGISTERS_15_22_port, B2 => n74, ZN => n884);
   U933 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n113_port, B1 => 
                           REGISTERS_11_22_port, B2 => n100_port, ZN => n883);
   U934 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n139, B1 => 
                           REGISTERS_14_22_port, B2 => n126_port, ZN => n882);
   U935 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n165, B1 => 
                           REGISTERS_10_22_port, B2 => n152, ZN => n881);
   U936 : NAND4_X1 port map( A1 => n884, A2 => n883, A3 => n882, A4 => n881, ZN
                           => n885);
   U937 : AOI22_X1 port map( A1 => n886, A2 => n1085, B1 => n885, B2 => n1083, 
                           ZN => n887);
   U938 : OAI221_X1 port map( B1 => n1089, B2 => n889, C1 => n1087, C2 => n888,
                           A => n887, ZN => N40);
   U939 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n87, B1 => 
                           REGISTERS_23_23_port, B2 => n74, ZN => n893);
   U940 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n113_port, B1 =>
                           REGISTERS_19_23_port, B2 => n100_port, ZN => n892);
   U941 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n139, B1 => 
                           REGISTERS_22_23_port, B2 => n126_port, ZN => n891);
   U942 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n165, B1 => 
                           REGISTERS_18_23_port, B2 => n152, ZN => n890);
   U943 : AND4_X1 port map( A1 => n893, A2 => n892, A3 => n891, A4 => n890, ZN 
                           => n910);
   U944 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n87, B1 => 
                           REGISTERS_31_23_port, B2 => n74, ZN => n897);
   U945 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n113_port, B1 =>
                           REGISTERS_27_23_port, B2 => n100_port, ZN => n896);
   U946 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n139, B1 => 
                           REGISTERS_30_23_port, B2 => n126_port, ZN => n895);
   U947 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n165, B1 => 
                           REGISTERS_26_23_port, B2 => n152, ZN => n894);
   U948 : AND4_X1 port map( A1 => n897, A2 => n896, A3 => n895, A4 => n894, ZN 
                           => n909);
   U949 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n87, B1 => 
                           REGISTERS_7_23_port, B2 => n74, ZN => n901);
   U950 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n113_port, B1 => 
                           REGISTERS_3_23_port, B2 => n100_port, ZN => n900);
   U951 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n139, B1 => 
                           REGISTERS_6_23_port, B2 => n126_port, ZN => n899);
   U952 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n165, B1 => 
                           REGISTERS_2_23_port, B2 => n152, ZN => n898);
   U953 : NAND4_X1 port map( A1 => n901, A2 => n900, A3 => n899, A4 => n898, ZN
                           => n907);
   U954 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n87, B1 => 
                           REGISTERS_15_23_port, B2 => n74, ZN => n905);
   U955 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n113_port, B1 => 
                           REGISTERS_11_23_port, B2 => n100_port, ZN => n904);
   U956 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n139, B1 => 
                           REGISTERS_14_23_port, B2 => n126_port, ZN => n903);
   U957 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n165, B1 => 
                           REGISTERS_10_23_port, B2 => n152, ZN => n902);
   U958 : NAND4_X1 port map( A1 => n905, A2 => n904, A3 => n903, A4 => n902, ZN
                           => n906);
   U959 : AOI22_X1 port map( A1 => n907, A2 => n1085, B1 => n906, B2 => n1083, 
                           ZN => n908);
   U960 : OAI221_X1 port map( B1 => n1089, B2 => n910, C1 => n1087, C2 => n909,
                           A => n908, ZN => N39);
   U961 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n88, B1 => 
                           REGISTERS_23_24_port, B2 => n75, ZN => n914);
   U962 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n114_port, B1 =>
                           REGISTERS_19_24_port, B2 => n101_port, ZN => n913);
   U963 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n140, B1 => 
                           REGISTERS_22_24_port, B2 => n127_port, ZN => n912);
   U964 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n166, B1 => 
                           REGISTERS_18_24_port, B2 => n153, ZN => n911);
   U965 : AND4_X1 port map( A1 => n914, A2 => n913, A3 => n912, A4 => n911, ZN 
                           => n931);
   U966 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n88, B1 => 
                           REGISTERS_31_24_port, B2 => n75, ZN => n918);
   U967 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n114_port, B1 =>
                           REGISTERS_27_24_port, B2 => n101_port, ZN => n917);
   U968 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n140, B1 => 
                           REGISTERS_30_24_port, B2 => n127_port, ZN => n916);
   U969 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n166, B1 => 
                           REGISTERS_26_24_port, B2 => n153, ZN => n915);
   U970 : AND4_X1 port map( A1 => n918, A2 => n917, A3 => n916, A4 => n915, ZN 
                           => n930);
   U971 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n88, B1 => 
                           REGISTERS_7_24_port, B2 => n75, ZN => n922);
   U972 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n114_port, B1 => 
                           REGISTERS_3_24_port, B2 => n101_port, ZN => n921);
   U973 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n140, B1 => 
                           REGISTERS_6_24_port, B2 => n127_port, ZN => n920);
   U974 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n166, B1 => 
                           REGISTERS_2_24_port, B2 => n153, ZN => n919);
   U975 : NAND4_X1 port map( A1 => n922, A2 => n921, A3 => n920, A4 => n919, ZN
                           => n928);
   U976 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n88, B1 => 
                           REGISTERS_15_24_port, B2 => n75, ZN => n926);
   U977 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n114_port, B1 => 
                           REGISTERS_11_24_port, B2 => n101_port, ZN => n925);
   U978 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n140, B1 => 
                           REGISTERS_14_24_port, B2 => n127_port, ZN => n924);
   U979 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n166, B1 => 
                           REGISTERS_10_24_port, B2 => n153, ZN => n923);
   U980 : NAND4_X1 port map( A1 => n926, A2 => n925, A3 => n924, A4 => n923, ZN
                           => n927);
   U981 : AOI22_X1 port map( A1 => n928, A2 => n1085, B1 => n927, B2 => n1083, 
                           ZN => n929);
   U982 : OAI221_X1 port map( B1 => n1089, B2 => n931, C1 => n1087, C2 => n930,
                           A => n929, ZN => N38);
   U983 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n88, B1 => 
                           REGISTERS_23_25_port, B2 => n75, ZN => n935);
   U984 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n114_port, B1 =>
                           REGISTERS_19_25_port, B2 => n101_port, ZN => n934);
   U985 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n140, B1 => 
                           REGISTERS_22_25_port, B2 => n127_port, ZN => n933);
   U986 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n166, B1 => 
                           REGISTERS_18_25_port, B2 => n153, ZN => n932);
   U987 : AND4_X1 port map( A1 => n935, A2 => n934, A3 => n933, A4 => n932, ZN 
                           => n952);
   U988 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n88, B1 => 
                           REGISTERS_31_25_port, B2 => n75, ZN => n939);
   U989 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n114_port, B1 =>
                           REGISTERS_27_25_port, B2 => n101_port, ZN => n938);
   U990 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n140, B1 => 
                           REGISTERS_30_25_port, B2 => n127_port, ZN => n937);
   U991 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n166, B1 => 
                           REGISTERS_26_25_port, B2 => n153, ZN => n936);
   U992 : AND4_X1 port map( A1 => n939, A2 => n938, A3 => n937, A4 => n936, ZN 
                           => n951);
   U993 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n88, B1 => 
                           REGISTERS_7_25_port, B2 => n75, ZN => n943);
   U994 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n114_port, B1 => 
                           REGISTERS_3_25_port, B2 => n101_port, ZN => n942);
   U995 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n140, B1 => 
                           REGISTERS_6_25_port, B2 => n127_port, ZN => n941);
   U996 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n166, B1 => 
                           REGISTERS_2_25_port, B2 => n153, ZN => n940);
   U997 : NAND4_X1 port map( A1 => n943, A2 => n942, A3 => n941, A4 => n940, ZN
                           => n949);
   U998 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n88, B1 => 
                           REGISTERS_15_25_port, B2 => n75, ZN => n947);
   U999 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n114_port, B1 => 
                           REGISTERS_11_25_port, B2 => n101_port, ZN => n946);
   U1000 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n140, B1 => 
                           REGISTERS_14_25_port, B2 => n127_port, ZN => n945);
   U1001 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n166, B1 => 
                           REGISTERS_10_25_port, B2 => n153, ZN => n944);
   U1002 : NAND4_X1 port map( A1 => n947, A2 => n946, A3 => n945, A4 => n944, 
                           ZN => n948);
   U1003 : AOI22_X1 port map( A1 => n949, A2 => n1085, B1 => n948, B2 => n1083,
                           ZN => n950);
   U1004 : OAI221_X1 port map( B1 => n1089, B2 => n952, C1 => n1087, C2 => n951
                           , A => n950, ZN => N37);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n88, B1 => 
                           REGISTERS_23_26_port, B2 => n75, ZN => n956);
   U1006 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n114_port, B1 
                           => REGISTERS_19_26_port, B2 => n101_port, ZN => n955
                           );
   U1007 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n140, B1 => 
                           REGISTERS_22_26_port, B2 => n127_port, ZN => n954);
   U1008 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n166, B1 => 
                           REGISTERS_18_26_port, B2 => n153, ZN => n953);
   U1009 : AND4_X1 port map( A1 => n956, A2 => n955, A3 => n954, A4 => n953, ZN
                           => n973);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n88, B1 => 
                           REGISTERS_31_26_port, B2 => n75, ZN => n960);
   U1011 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n114_port, B1 
                           => REGISTERS_27_26_port, B2 => n101_port, ZN => n959
                           );
   U1012 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n140, B1 => 
                           REGISTERS_30_26_port, B2 => n127_port, ZN => n958);
   U1013 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n166, B1 => 
                           REGISTERS_26_26_port, B2 => n153, ZN => n957);
   U1014 : AND4_X1 port map( A1 => n960, A2 => n959, A3 => n958, A4 => n957, ZN
                           => n972);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n88, B1 => 
                           REGISTERS_7_26_port, B2 => n75, ZN => n964);
   U1016 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n114_port, B1 =>
                           REGISTERS_3_26_port, B2 => n101_port, ZN => n963);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n140, B1 => 
                           REGISTERS_6_26_port, B2 => n127_port, ZN => n962);
   U1018 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n166, B1 => 
                           REGISTERS_2_26_port, B2 => n153, ZN => n961);
   U1019 : NAND4_X1 port map( A1 => n964, A2 => n963, A3 => n962, A4 => n961, 
                           ZN => n970);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n88, B1 => 
                           REGISTERS_15_26_port, B2 => n75, ZN => n968);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n114_port, B1 =>
                           REGISTERS_11_26_port, B2 => n101_port, ZN => n967);
   U1022 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n140, B1 => 
                           REGISTERS_14_26_port, B2 => n127_port, ZN => n966);
   U1023 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n166, B1 => 
                           REGISTERS_10_26_port, B2 => n153, ZN => n965);
   U1024 : NAND4_X1 port map( A1 => n968, A2 => n967, A3 => n966, A4 => n965, 
                           ZN => n969);
   U1025 : AOI22_X1 port map( A1 => n970, A2 => n1085, B1 => n969, B2 => n1083,
                           ZN => n971);
   U1026 : OAI221_X1 port map( B1 => n1089, B2 => n973, C1 => n1087, C2 => n972
                           , A => n971, ZN => N36);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n89, B1 => 
                           REGISTERS_23_27_port, B2 => n76, ZN => n977);
   U1028 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n115_port, B1 
                           => REGISTERS_19_27_port, B2 => n102_port, ZN => n976
                           );
   U1029 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n141, B1 => 
                           REGISTERS_22_27_port, B2 => n128, ZN => n975);
   U1030 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n167, B1 => 
                           REGISTERS_18_27_port, B2 => n154, ZN => n974);
   U1031 : AND4_X1 port map( A1 => n977, A2 => n976, A3 => n975, A4 => n974, ZN
                           => n994);
   U1032 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n89, B1 => 
                           REGISTERS_31_27_port, B2 => n76, ZN => n981);
   U1033 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n115_port, B1 
                           => REGISTERS_27_27_port, B2 => n102_port, ZN => n980
                           );
   U1034 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n141, B1 => 
                           REGISTERS_30_27_port, B2 => n128, ZN => n979);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n167, B1 => 
                           REGISTERS_26_27_port, B2 => n154, ZN => n978);
   U1036 : AND4_X1 port map( A1 => n981, A2 => n980, A3 => n979, A4 => n978, ZN
                           => n993);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n89, B1 => 
                           REGISTERS_7_27_port, B2 => n76, ZN => n985);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n115_port, B1 =>
                           REGISTERS_3_27_port, B2 => n102_port, ZN => n984);
   U1039 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n141, B1 => 
                           REGISTERS_6_27_port, B2 => n128, ZN => n983);
   U1040 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n167, B1 => 
                           REGISTERS_2_27_port, B2 => n154, ZN => n982);
   U1041 : NAND4_X1 port map( A1 => n985, A2 => n984, A3 => n983, A4 => n982, 
                           ZN => n991);
   U1042 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n89, B1 => 
                           REGISTERS_15_27_port, B2 => n76, ZN => n989);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n115_port, B1 =>
                           REGISTERS_11_27_port, B2 => n102_port, ZN => n988);
   U1044 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n141, B1 => 
                           REGISTERS_14_27_port, B2 => n128, ZN => n987);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n167, B1 => 
                           REGISTERS_10_27_port, B2 => n154, ZN => n986);
   U1046 : NAND4_X1 port map( A1 => n989, A2 => n988, A3 => n987, A4 => n986, 
                           ZN => n990);
   U1047 : AOI22_X1 port map( A1 => n991, A2 => n1085, B1 => n990, B2 => n1083,
                           ZN => n992);
   U1048 : OAI221_X1 port map( B1 => n1089, B2 => n994, C1 => n1087, C2 => n993
                           , A => n992, ZN => N35);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n89, B1 => 
                           REGISTERS_23_28_port, B2 => n76, ZN => n998);
   U1050 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n115_port, B1 
                           => REGISTERS_19_28_port, B2 => n102_port, ZN => n997
                           );
   U1051 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n141, B1 => 
                           REGISTERS_22_28_port, B2 => n128, ZN => n996);
   U1052 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n167, B1 => 
                           REGISTERS_18_28_port, B2 => n154, ZN => n995);
   U1053 : AND4_X1 port map( A1 => n998, A2 => n997, A3 => n996, A4 => n995, ZN
                           => n1015);
   U1054 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n89, B1 => 
                           REGISTERS_31_28_port, B2 => n76, ZN => n1002);
   U1055 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n115_port, B1 
                           => REGISTERS_27_28_port, B2 => n102_port, ZN => 
                           n1001);
   U1056 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n141, B1 => 
                           REGISTERS_30_28_port, B2 => n128, ZN => n1000);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n167, B1 => 
                           REGISTERS_26_28_port, B2 => n154, ZN => n999);
   U1058 : AND4_X1 port map( A1 => n1002, A2 => n1001, A3 => n1000, A4 => n999,
                           ZN => n1014);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n89, B1 => 
                           REGISTERS_7_28_port, B2 => n76, ZN => n1006);
   U1060 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n115_port, B1 =>
                           REGISTERS_3_28_port, B2 => n102_port, ZN => n1005);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n141, B1 => 
                           REGISTERS_6_28_port, B2 => n128, ZN => n1004);
   U1062 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n167, B1 => 
                           REGISTERS_2_28_port, B2 => n154, ZN => n1003);
   U1063 : NAND4_X1 port map( A1 => n1006, A2 => n1005, A3 => n1004, A4 => 
                           n1003, ZN => n1012);
   U1064 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n89, B1 => 
                           REGISTERS_15_28_port, B2 => n76, ZN => n1010);
   U1065 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n115_port, B1 =>
                           REGISTERS_11_28_port, B2 => n102_port, ZN => n1009);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n141, B1 => 
                           REGISTERS_14_28_port, B2 => n128, ZN => n1008);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n167, B1 => 
                           REGISTERS_10_28_port, B2 => n154, ZN => n1007);
   U1068 : NAND4_X1 port map( A1 => n1010, A2 => n1009, A3 => n1008, A4 => 
                           n1007, ZN => n1011);
   U1069 : AOI22_X1 port map( A1 => n1012, A2 => n1085, B1 => n1011, B2 => 
                           n1083, ZN => n1013);
   U1070 : OAI221_X1 port map( B1 => n1089, B2 => n1015, C1 => n1087, C2 => 
                           n1014, A => n1013, ZN => N34);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n89, B1 => 
                           REGISTERS_23_29_port, B2 => n76, ZN => n1019);
   U1072 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n115_port, B1 
                           => REGISTERS_19_29_port, B2 => n102_port, ZN => 
                           n1018);
   U1073 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n141, B1 => 
                           REGISTERS_22_29_port, B2 => n128, ZN => n1017);
   U1074 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n167, B1 => 
                           REGISTERS_18_29_port, B2 => n154, ZN => n1016);
   U1075 : AND4_X1 port map( A1 => n1019, A2 => n1018, A3 => n1017, A4 => n1016
                           , ZN => n1036);
   U1076 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n89, B1 => 
                           REGISTERS_31_29_port, B2 => n76, ZN => n1023);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n115_port, B1 
                           => REGISTERS_27_29_port, B2 => n102_port, ZN => 
                           n1022);
   U1078 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n141, B1 => 
                           REGISTERS_30_29_port, B2 => n128, ZN => n1021);
   U1079 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n167, B1 => 
                           REGISTERS_26_29_port, B2 => n154, ZN => n1020);
   U1080 : AND4_X1 port map( A1 => n1023, A2 => n1022, A3 => n1021, A4 => n1020
                           , ZN => n1035);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n89, B1 => 
                           REGISTERS_7_29_port, B2 => n76, ZN => n1027);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n115_port, B1 =>
                           REGISTERS_3_29_port, B2 => n102_port, ZN => n1026);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n141, B1 => 
                           REGISTERS_6_29_port, B2 => n128, ZN => n1025);
   U1084 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n167, B1 => 
                           REGISTERS_2_29_port, B2 => n154, ZN => n1024);
   U1085 : NAND4_X1 port map( A1 => n1027, A2 => n1026, A3 => n1025, A4 => 
                           n1024, ZN => n1033);
   U1086 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n89, B1 => 
                           REGISTERS_15_29_port, B2 => n76, ZN => n1031);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n115_port, B1 =>
                           REGISTERS_11_29_port, B2 => n102_port, ZN => n1030);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n141, B1 => 
                           REGISTERS_14_29_port, B2 => n128, ZN => n1029);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n167, B1 => 
                           REGISTERS_10_29_port, B2 => n154, ZN => n1028);
   U1090 : NAND4_X1 port map( A1 => n1031, A2 => n1030, A3 => n1029, A4 => 
                           n1028, ZN => n1032);
   U1091 : AOI22_X1 port map( A1 => n1033, A2 => n1085, B1 => n1032, B2 => 
                           n1083, ZN => n1034);
   U1092 : OAI221_X1 port map( B1 => n1089, B2 => n1036, C1 => n1087, C2 => 
                           n1035, A => n1034, ZN => N33);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n90, B1 => 
                           REGISTERS_23_30_port, B2 => n77, ZN => n1040);
   U1094 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n116_port, B1 
                           => REGISTERS_19_30_port, B2 => n103_port, ZN => 
                           n1039);
   U1095 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n142, B1 => 
                           REGISTERS_22_30_port, B2 => n129, ZN => n1038);
   U1096 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n168, B1 => 
                           REGISTERS_18_30_port, B2 => n155, ZN => n1037);
   U1097 : AND4_X1 port map( A1 => n1040, A2 => n1039, A3 => n1038, A4 => n1037
                           , ZN => n1057);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n90, B1 => 
                           REGISTERS_31_30_port, B2 => n77, ZN => n1044);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n116_port, B1 
                           => REGISTERS_27_30_port, B2 => n103_port, ZN => 
                           n1043);
   U1100 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n142, B1 => 
                           REGISTERS_30_30_port, B2 => n129, ZN => n1042);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n168, B1 => 
                           REGISTERS_26_30_port, B2 => n155, ZN => n1041);
   U1102 : AND4_X1 port map( A1 => n1044, A2 => n1043, A3 => n1042, A4 => n1041
                           , ZN => n1056);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n90, B1 => 
                           REGISTERS_7_30_port, B2 => n77, ZN => n1048);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n116_port, B1 =>
                           REGISTERS_3_30_port, B2 => n103_port, ZN => n1047);
   U1105 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n142, B1 => 
                           REGISTERS_6_30_port, B2 => n129, ZN => n1046);
   U1106 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n168, B1 => 
                           REGISTERS_2_30_port, B2 => n155, ZN => n1045);
   U1107 : NAND4_X1 port map( A1 => n1048, A2 => n1047, A3 => n1046, A4 => 
                           n1045, ZN => n1054);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n90, B1 => 
                           REGISTERS_15_30_port, B2 => n77, ZN => n1052);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n116_port, B1 =>
                           REGISTERS_11_30_port, B2 => n103_port, ZN => n1051);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n142, B1 => 
                           REGISTERS_14_30_port, B2 => n129, ZN => n1050);
   U1111 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n168, B1 => 
                           REGISTERS_10_30_port, B2 => n155, ZN => n1049);
   U1112 : NAND4_X1 port map( A1 => n1052, A2 => n1051, A3 => n1050, A4 => 
                           n1049, ZN => n1053);
   U1113 : AOI22_X1 port map( A1 => n1054, A2 => n1085, B1 => n1053, B2 => 
                           n1083, ZN => n1055);
   U1114 : OAI221_X1 port map( B1 => n1089, B2 => n1057, C1 => n1087, C2 => 
                           n1056, A => n1055, ZN => N32);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n90, B1 => 
                           REGISTERS_23_31_port, B2 => n77, ZN => n1061);
   U1116 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n116_port, B1 
                           => REGISTERS_19_31_port, B2 => n103_port, ZN => 
                           n1060);
   U1117 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n142, B1 => 
                           REGISTERS_22_31_port, B2 => n129, ZN => n1059);
   U1118 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n168, B1 => 
                           REGISTERS_18_31_port, B2 => n155, ZN => n1058);
   U1119 : AND4_X1 port map( A1 => n1061, A2 => n1060, A3 => n1059, A4 => n1058
                           , ZN => n1090);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n90, B1 => 
                           REGISTERS_31_31_port, B2 => n77, ZN => n1065);
   U1121 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n116_port, B1 
                           => REGISTERS_27_31_port, B2 => n103_port, ZN => 
                           n1064);
   U1122 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n142, B1 => 
                           REGISTERS_30_31_port, B2 => n129, ZN => n1063);
   U1123 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n168, B1 => 
                           REGISTERS_26_31_port, B2 => n155, ZN => n1062);
   U1124 : AND4_X1 port map( A1 => n1065, A2 => n1064, A3 => n1063, A4 => n1062
                           , ZN => n1088);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n90, B1 => 
                           REGISTERS_7_31_port, B2 => n77, ZN => n1069);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n116_port, B1 =>
                           REGISTERS_3_31_port, B2 => n103_port, ZN => n1068);
   U1127 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n142, B1 => 
                           REGISTERS_6_31_port, B2 => n129, ZN => n1067);
   U1128 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n168, B1 => 
                           REGISTERS_2_31_port, B2 => n155, ZN => n1066);
   U1129 : NAND4_X1 port map( A1 => n1069, A2 => n1068, A3 => n1067, A4 => 
                           n1066, ZN => n1084);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n90, B1 => 
                           REGISTERS_15_31_port, B2 => n77, ZN => n1081);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n116_port, B1 =>
                           REGISTERS_11_31_port, B2 => n103_port, ZN => n1080);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n142, B1 => 
                           REGISTERS_14_31_port, B2 => n129, ZN => n1079);
   U1133 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n168, B1 => 
                           REGISTERS_10_31_port, B2 => n155, ZN => n1078);
   U1134 : NAND4_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, A4 => 
                           n1078, ZN => n1082);
   U1135 : AOI22_X1 port map( A1 => n1085, A2 => n1084, B1 => n1083, B2 => 
                           n1082, ZN => n1086);
   U1136 : OAI221_X1 port map( B1 => n1090, B2 => n1089, C1 => n1088, C2 => 
                           n1087, A => n1086, ZN => N31);
   U1137 : NOR2_X1 port map( A1 => n2808, A2 => ADD_RD2(1), ZN => n1095);
   U1138 : AND2_X1 port map( A1 => n1095, A2 => ADD_RD2(0), ZN => n2787);
   U1139 : NOR2_X1 port map( A1 => n2808, A2 => n2809, ZN => n1096);
   U1140 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1096, ZN => n2786);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n184, B1 => 
                           REGISTERS_23_0_port, B2 => n171, ZN => n1102);
   U1142 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1097);
   U1143 : AND2_X1 port map( A1 => n1097, A2 => ADD_RD2(0), ZN => n2789);
   U1144 : NOR2_X1 port map( A1 => n2809, A2 => ADD_RD2(2), ZN => n1098);
   U1145 : AND2_X1 port map( A1 => n1098, A2 => ADD_RD2(0), ZN => n2788);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n210, B1 => 
                           REGISTERS_19_0_port, B2 => n197, ZN => n1101);
   U1147 : AND2_X1 port map( A1 => n1095, A2 => n2810, ZN => n2791);
   U1148 : AND2_X1 port map( A1 => n1096, A2 => n2810, ZN => n2790);
   U1149 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n236, B1 => 
                           REGISTERS_22_0_port, B2 => n223, ZN => n1100);
   U1150 : AND2_X1 port map( A1 => n1097, A2 => n2810, ZN => n2793);
   U1151 : AND2_X1 port map( A1 => n1098, A2 => n2810, ZN => n2792);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n262, B1 => 
                           REGISTERS_18_0_port, B2 => n249, ZN => n1099);
   U1153 : AND4_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, A4 => n1099
                           , ZN => n1119);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n184, B1 => 
                           REGISTERS_31_0_port, B2 => n171, ZN => n1106);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n210, B1 => 
                           REGISTERS_27_0_port, B2 => n197, ZN => n1105);
   U1156 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n236, B1 => 
                           REGISTERS_30_0_port, B2 => n223, ZN => n1104);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n262, B1 => 
                           REGISTERS_26_0_port, B2 => n249, ZN => n1103);
   U1158 : AND4_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, A4 => n1103
                           , ZN => n1118);
   U1159 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n184, B1 => 
                           REGISTERS_7_0_port, B2 => n171, ZN => n1110);
   U1160 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n210, B1 => 
                           REGISTERS_3_0_port, B2 => n197, ZN => n1109);
   U1161 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n236, B1 => 
                           REGISTERS_6_0_port, B2 => n223, ZN => n1108);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n262, B1 => 
                           REGISTERS_2_0_port, B2 => n249, ZN => n1107);
   U1163 : NAND4_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, A4 => 
                           n1107, ZN => n1116);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n184, B1 => 
                           REGISTERS_15_0_port, B2 => n171, ZN => n1114);
   U1165 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n210, B1 => 
                           REGISTERS_11_0_port, B2 => n197, ZN => n1113);
   U1166 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n236, B1 => 
                           REGISTERS_14_0_port, B2 => n223, ZN => n1112);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n262, B1 => 
                           REGISTERS_10_0_port, B2 => n249, ZN => n1111);
   U1168 : NAND4_X1 port map( A1 => n1114, A2 => n1113, A3 => n1112, A4 => 
                           n1111, ZN => n1115);
   U1169 : AOI22_X1 port map( A1 => n1116, A2 => n2801, B1 => n1115, B2 => 
                           n2799, ZN => n1117);
   U1170 : OAI221_X1 port map( B1 => n2805, B2 => n1119, C1 => n2803, C2 => 
                           n1118, A => n1117, ZN => N127);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n184, B1 => 
                           REGISTERS_23_1_port, B2 => n171, ZN => n1123);
   U1172 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n210, B1 => 
                           REGISTERS_19_1_port, B2 => n197, ZN => n1122);
   U1173 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n236, B1 => 
                           REGISTERS_22_1_port, B2 => n223, ZN => n1121);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n262, B1 => 
                           REGISTERS_18_1_port, B2 => n249, ZN => n1120);
   U1175 : AND4_X1 port map( A1 => n1123, A2 => n1122, A3 => n1121, A4 => n1120
                           , ZN => n1140);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n184, B1 => 
                           REGISTERS_31_1_port, B2 => n171, ZN => n1127);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n210, B1 => 
                           REGISTERS_27_1_port, B2 => n197, ZN => n1126);
   U1178 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n236, B1 => 
                           REGISTERS_30_1_port, B2 => n223, ZN => n1125);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n262, B1 => 
                           REGISTERS_26_1_port, B2 => n249, ZN => n1124);
   U1180 : AND4_X1 port map( A1 => n1127, A2 => n1126, A3 => n1125, A4 => n1124
                           , ZN => n1139);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n184, B1 => 
                           REGISTERS_7_1_port, B2 => n171, ZN => n1131);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n210, B1 => 
                           REGISTERS_3_1_port, B2 => n197, ZN => n1130);
   U1183 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n236, B1 => 
                           REGISTERS_6_1_port, B2 => n223, ZN => n1129);
   U1184 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n262, B1 => 
                           REGISTERS_2_1_port, B2 => n249, ZN => n1128);
   U1185 : NAND4_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, A4 => 
                           n1128, ZN => n1137);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n184, B1 => 
                           REGISTERS_15_1_port, B2 => n171, ZN => n1135);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n210, B1 => 
                           REGISTERS_11_1_port, B2 => n197, ZN => n1134);
   U1188 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n236, B1 => 
                           REGISTERS_14_1_port, B2 => n223, ZN => n1133);
   U1189 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n262, B1 => 
                           REGISTERS_10_1_port, B2 => n249, ZN => n1132);
   U1190 : NAND4_X1 port map( A1 => n1135, A2 => n1134, A3 => n1133, A4 => 
                           n1132, ZN => n1136);
   U1191 : AOI22_X1 port map( A1 => n1137, A2 => n2801, B1 => n1136, B2 => 
                           n2799, ZN => n1138);
   U1192 : OAI221_X1 port map( B1 => n2805, B2 => n1140, C1 => n2803, C2 => 
                           n1139, A => n1138, ZN => N126);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n184, B1 => 
                           REGISTERS_23_2_port, B2 => n171, ZN => n2168);
   U1194 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n210, B1 => 
                           REGISTERS_19_2_port, B2 => n197, ZN => n2167);
   U1195 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n236, B1 => 
                           REGISTERS_22_2_port, B2 => n223, ZN => n1142);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n262, B1 => 
                           REGISTERS_18_2_port, B2 => n249, ZN => n1141);
   U1197 : AND4_X1 port map( A1 => n2168, A2 => n2167, A3 => n1142, A4 => n1141
                           , ZN => n2185);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n184, B1 => 
                           REGISTERS_31_2_port, B2 => n171, ZN => n2172);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n210, B1 => 
                           REGISTERS_27_2_port, B2 => n197, ZN => n2171);
   U1200 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n236, B1 => 
                           REGISTERS_30_2_port, B2 => n223, ZN => n2170);
   U1201 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n262, B1 => 
                           REGISTERS_26_2_port, B2 => n249, ZN => n2169);
   U1202 : AND4_X1 port map( A1 => n2172, A2 => n2171, A3 => n2170, A4 => n2169
                           , ZN => n2184);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n184, B1 => 
                           REGISTERS_7_2_port, B2 => n171, ZN => n2176);
   U1204 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n210, B1 => 
                           REGISTERS_3_2_port, B2 => n197, ZN => n2175);
   U1205 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n236, B1 => 
                           REGISTERS_6_2_port, B2 => n223, ZN => n2174);
   U1206 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n262, B1 => 
                           REGISTERS_2_2_port, B2 => n249, ZN => n2173);
   U1207 : NAND4_X1 port map( A1 => n2176, A2 => n2175, A3 => n2174, A4 => 
                           n2173, ZN => n2182);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n184, B1 => 
                           REGISTERS_15_2_port, B2 => n171, ZN => n2180);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n210, B1 => 
                           REGISTERS_11_2_port, B2 => n197, ZN => n2179);
   U1210 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n236, B1 => 
                           REGISTERS_14_2_port, B2 => n223, ZN => n2178);
   U1211 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n262, B1 => 
                           REGISTERS_10_2_port, B2 => n249, ZN => n2177);
   U1212 : NAND4_X1 port map( A1 => n2180, A2 => n2179, A3 => n2178, A4 => 
                           n2177, ZN => n2181);
   U1213 : AOI22_X1 port map( A1 => n2182, A2 => n2801, B1 => n2181, B2 => 
                           n2799, ZN => n2183);
   U1214 : OAI221_X1 port map( B1 => n2805, B2 => n2185, C1 => n2803, C2 => 
                           n2184, A => n2183, ZN => N125);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n185, B1 => 
                           REGISTERS_23_3_port, B2 => n172, ZN => n2189);
   U1216 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n211, B1 => 
                           REGISTERS_19_3_port, B2 => n198, ZN => n2188);
   U1217 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n237, B1 => 
                           REGISTERS_22_3_port, B2 => n224, ZN => n2187);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n263, B1 => 
                           REGISTERS_18_3_port, B2 => n250, ZN => n2186);
   U1219 : AND4_X1 port map( A1 => n2189, A2 => n2188, A3 => n2187, A4 => n2186
                           , ZN => n2206);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n185, B1 => 
                           REGISTERS_31_3_port, B2 => n172, ZN => n2193);
   U1221 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n211, B1 => 
                           REGISTERS_27_3_port, B2 => n198, ZN => n2192);
   U1222 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n237, B1 => 
                           REGISTERS_30_3_port, B2 => n224, ZN => n2191);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n263, B1 => 
                           REGISTERS_26_3_port, B2 => n250, ZN => n2190);
   U1224 : AND4_X1 port map( A1 => n2193, A2 => n2192, A3 => n2191, A4 => n2190
                           , ZN => n2205);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n185, B1 => 
                           REGISTERS_7_3_port, B2 => n172, ZN => n2197);
   U1226 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n211, B1 => 
                           REGISTERS_3_3_port, B2 => n198, ZN => n2196);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n237, B1 => 
                           REGISTERS_6_3_port, B2 => n224, ZN => n2195);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n263, B1 => 
                           REGISTERS_2_3_port, B2 => n250, ZN => n2194);
   U1229 : NAND4_X1 port map( A1 => n2197, A2 => n2196, A3 => n2195, A4 => 
                           n2194, ZN => n2203);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n185, B1 => 
                           REGISTERS_15_3_port, B2 => n172, ZN => n2201);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n211, B1 => 
                           REGISTERS_11_3_port, B2 => n198, ZN => n2200);
   U1232 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n237, B1 => 
                           REGISTERS_14_3_port, B2 => n224, ZN => n2199);
   U1233 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n263, B1 => 
                           REGISTERS_10_3_port, B2 => n250, ZN => n2198);
   U1234 : NAND4_X1 port map( A1 => n2201, A2 => n2200, A3 => n2199, A4 => 
                           n2198, ZN => n2202);
   U1235 : AOI22_X1 port map( A1 => n2203, A2 => n2801, B1 => n2202, B2 => 
                           n2799, ZN => n2204);
   U1236 : OAI221_X1 port map( B1 => n2805, B2 => n2206, C1 => n2803, C2 => 
                           n2205, A => n2204, ZN => N124);
   U1237 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n185, B1 => 
                           REGISTERS_23_4_port, B2 => n172, ZN => n2210);
   U1238 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n211, B1 => 
                           REGISTERS_19_4_port, B2 => n198, ZN => n2209);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n237, B1 => 
                           REGISTERS_22_4_port, B2 => n224, ZN => n2208);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n263, B1 => 
                           REGISTERS_18_4_port, B2 => n250, ZN => n2207);
   U1241 : AND4_X1 port map( A1 => n2210, A2 => n2209, A3 => n2208, A4 => n2207
                           , ZN => n2227);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n185, B1 => 
                           REGISTERS_31_4_port, B2 => n172, ZN => n2214);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n211, B1 => 
                           REGISTERS_27_4_port, B2 => n198, ZN => n2213);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n237, B1 => 
                           REGISTERS_30_4_port, B2 => n224, ZN => n2212);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n263, B1 => 
                           REGISTERS_26_4_port, B2 => n250, ZN => n2211);
   U1246 : AND4_X1 port map( A1 => n2214, A2 => n2213, A3 => n2212, A4 => n2211
                           , ZN => n2226);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n185, B1 => 
                           REGISTERS_7_4_port, B2 => n172, ZN => n2218);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n211, B1 => 
                           REGISTERS_3_4_port, B2 => n198, ZN => n2217);
   U1249 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n237, B1 => 
                           REGISTERS_6_4_port, B2 => n224, ZN => n2216);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n263, B1 => 
                           REGISTERS_2_4_port, B2 => n250, ZN => n2215);
   U1251 : NAND4_X1 port map( A1 => n2218, A2 => n2217, A3 => n2216, A4 => 
                           n2215, ZN => n2224);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n185, B1 => 
                           REGISTERS_15_4_port, B2 => n172, ZN => n2222);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n211, B1 => 
                           REGISTERS_11_4_port, B2 => n198, ZN => n2221);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n237, B1 => 
                           REGISTERS_14_4_port, B2 => n224, ZN => n2220);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n263, B1 => 
                           REGISTERS_10_4_port, B2 => n250, ZN => n2219);
   U1256 : NAND4_X1 port map( A1 => n2222, A2 => n2221, A3 => n2220, A4 => 
                           n2219, ZN => n2223);
   U1257 : AOI22_X1 port map( A1 => n2224, A2 => n2801, B1 => n2223, B2 => 
                           n2799, ZN => n2225);
   U1258 : OAI221_X1 port map( B1 => n2805, B2 => n2227, C1 => n2803, C2 => 
                           n2226, A => n2225, ZN => N123);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n185, B1 => 
                           REGISTERS_23_5_port, B2 => n172, ZN => n2231);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n211, B1 => 
                           REGISTERS_19_5_port, B2 => n198, ZN => n2230);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n237, B1 => 
                           REGISTERS_22_5_port, B2 => n224, ZN => n2229);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n263, B1 => 
                           REGISTERS_18_5_port, B2 => n250, ZN => n2228);
   U1263 : AND4_X1 port map( A1 => n2231, A2 => n2230, A3 => n2229, A4 => n2228
                           , ZN => n2248);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n185, B1 => 
                           REGISTERS_31_5_port, B2 => n172, ZN => n2235);
   U1265 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n211, B1 => 
                           REGISTERS_27_5_port, B2 => n198, ZN => n2234);
   U1266 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n237, B1 => 
                           REGISTERS_30_5_port, B2 => n224, ZN => n2233);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n263, B1 => 
                           REGISTERS_26_5_port, B2 => n250, ZN => n2232);
   U1268 : AND4_X1 port map( A1 => n2235, A2 => n2234, A3 => n2233, A4 => n2232
                           , ZN => n2247);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n185, B1 => 
                           REGISTERS_7_5_port, B2 => n172, ZN => n2239);
   U1270 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n211, B1 => 
                           REGISTERS_3_5_port, B2 => n198, ZN => n2238);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n237, B1 => 
                           REGISTERS_6_5_port, B2 => n224, ZN => n2237);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n263, B1 => 
                           REGISTERS_2_5_port, B2 => n250, ZN => n2236);
   U1273 : NAND4_X1 port map( A1 => n2239, A2 => n2238, A3 => n2237, A4 => 
                           n2236, ZN => n2245);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n185, B1 => 
                           REGISTERS_15_5_port, B2 => n172, ZN => n2243);
   U1275 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n211, B1 => 
                           REGISTERS_11_5_port, B2 => n198, ZN => n2242);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n237, B1 => 
                           REGISTERS_14_5_port, B2 => n224, ZN => n2241);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n263, B1 => 
                           REGISTERS_10_5_port, B2 => n250, ZN => n2240);
   U1278 : NAND4_X1 port map( A1 => n2243, A2 => n2242, A3 => n2241, A4 => 
                           n2240, ZN => n2244);
   U1279 : AOI22_X1 port map( A1 => n2245, A2 => n2801, B1 => n2244, B2 => 
                           n2799, ZN => n2246);
   U1280 : OAI221_X1 port map( B1 => n2805, B2 => n2248, C1 => n2803, C2 => 
                           n2247, A => n2246, ZN => N122);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n186, B1 => 
                           REGISTERS_23_6_port, B2 => n173, ZN => n2252);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n212, B1 => 
                           REGISTERS_19_6_port, B2 => n199, ZN => n2251);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n238, B1 => 
                           REGISTERS_22_6_port, B2 => n225, ZN => n2250);
   U1284 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n264, B1 => 
                           REGISTERS_18_6_port, B2 => n251, ZN => n2249);
   U1285 : AND4_X1 port map( A1 => n2252, A2 => n2251, A3 => n2250, A4 => n2249
                           , ZN => n2269);
   U1286 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n186, B1 => 
                           REGISTERS_31_6_port, B2 => n173, ZN => n2256);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n212, B1 => 
                           REGISTERS_27_6_port, B2 => n199, ZN => n2255);
   U1288 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n238, B1 => 
                           REGISTERS_30_6_port, B2 => n225, ZN => n2254);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n264, B1 => 
                           REGISTERS_26_6_port, B2 => n251, ZN => n2253);
   U1290 : AND4_X1 port map( A1 => n2256, A2 => n2255, A3 => n2254, A4 => n2253
                           , ZN => n2268);
   U1291 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n186, B1 => 
                           REGISTERS_7_6_port, B2 => n173, ZN => n2260);
   U1292 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n212, B1 => 
                           REGISTERS_3_6_port, B2 => n199, ZN => n2259);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n238, B1 => 
                           REGISTERS_6_6_port, B2 => n225, ZN => n2258);
   U1294 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n264, B1 => 
                           REGISTERS_2_6_port, B2 => n251, ZN => n2257);
   U1295 : NAND4_X1 port map( A1 => n2260, A2 => n2259, A3 => n2258, A4 => 
                           n2257, ZN => n2266);
   U1296 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n186, B1 => 
                           REGISTERS_15_6_port, B2 => n173, ZN => n2264);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n212, B1 => 
                           REGISTERS_11_6_port, B2 => n199, ZN => n2263);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n238, B1 => 
                           REGISTERS_14_6_port, B2 => n225, ZN => n2262);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n264, B1 => 
                           REGISTERS_10_6_port, B2 => n251, ZN => n2261);
   U1300 : NAND4_X1 port map( A1 => n2264, A2 => n2263, A3 => n2262, A4 => 
                           n2261, ZN => n2265);
   U1301 : AOI22_X1 port map( A1 => n2266, A2 => n2801, B1 => n2265, B2 => 
                           n2799, ZN => n2267);
   U1302 : OAI221_X1 port map( B1 => n2805, B2 => n2269, C1 => n2803, C2 => 
                           n2268, A => n2267, ZN => N121);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n186, B1 => 
                           REGISTERS_23_7_port, B2 => n173, ZN => n2273);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n212, B1 => 
                           REGISTERS_19_7_port, B2 => n199, ZN => n2272);
   U1305 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n238, B1 => 
                           REGISTERS_22_7_port, B2 => n225, ZN => n2271);
   U1306 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n264, B1 => 
                           REGISTERS_18_7_port, B2 => n251, ZN => n2270);
   U1307 : AND4_X1 port map( A1 => n2273, A2 => n2272, A3 => n2271, A4 => n2270
                           , ZN => n2290);
   U1308 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n186, B1 => 
                           REGISTERS_31_7_port, B2 => n173, ZN => n2277);
   U1309 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n212, B1 => 
                           REGISTERS_27_7_port, B2 => n199, ZN => n2276);
   U1310 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n238, B1 => 
                           REGISTERS_30_7_port, B2 => n225, ZN => n2275);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n264, B1 => 
                           REGISTERS_26_7_port, B2 => n251, ZN => n2274);
   U1312 : AND4_X1 port map( A1 => n2277, A2 => n2276, A3 => n2275, A4 => n2274
                           , ZN => n2289);
   U1313 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n186, B1 => 
                           REGISTERS_7_7_port, B2 => n173, ZN => n2281);
   U1314 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n212, B1 => 
                           REGISTERS_3_7_port, B2 => n199, ZN => n2280);
   U1315 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n238, B1 => 
                           REGISTERS_6_7_port, B2 => n225, ZN => n2279);
   U1316 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n264, B1 => 
                           REGISTERS_2_7_port, B2 => n251, ZN => n2278);
   U1317 : NAND4_X1 port map( A1 => n2281, A2 => n2280, A3 => n2279, A4 => 
                           n2278, ZN => n2287);
   U1318 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n186, B1 => 
                           REGISTERS_15_7_port, B2 => n173, ZN => n2285);
   U1319 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n212, B1 => 
                           REGISTERS_11_7_port, B2 => n199, ZN => n2284);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n238, B1 => 
                           REGISTERS_14_7_port, B2 => n225, ZN => n2283);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n264, B1 => 
                           REGISTERS_10_7_port, B2 => n251, ZN => n2282);
   U1322 : NAND4_X1 port map( A1 => n2285, A2 => n2284, A3 => n2283, A4 => 
                           n2282, ZN => n2286);
   U1323 : AOI22_X1 port map( A1 => n2287, A2 => n2801, B1 => n2286, B2 => 
                           n2799, ZN => n2288);
   U1324 : OAI221_X1 port map( B1 => n2805, B2 => n2290, C1 => n2803, C2 => 
                           n2289, A => n2288, ZN => N120);
   U1325 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n186, B1 => 
                           REGISTERS_23_8_port, B2 => n173, ZN => n2294);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n212, B1 => 
                           REGISTERS_19_8_port, B2 => n199, ZN => n2293);
   U1327 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n238, B1 => 
                           REGISTERS_22_8_port, B2 => n225, ZN => n2292);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n264, B1 => 
                           REGISTERS_18_8_port, B2 => n251, ZN => n2291);
   U1329 : AND4_X1 port map( A1 => n2294, A2 => n2293, A3 => n2292, A4 => n2291
                           , ZN => n2311);
   U1330 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n186, B1 => 
                           REGISTERS_31_8_port, B2 => n173, ZN => n2298);
   U1331 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n212, B1 => 
                           REGISTERS_27_8_port, B2 => n199, ZN => n2297);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n238, B1 => 
                           REGISTERS_30_8_port, B2 => n225, ZN => n2296);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n264, B1 => 
                           REGISTERS_26_8_port, B2 => n251, ZN => n2295);
   U1334 : AND4_X1 port map( A1 => n2298, A2 => n2297, A3 => n2296, A4 => n2295
                           , ZN => n2310);
   U1335 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n186, B1 => 
                           REGISTERS_7_8_port, B2 => n173, ZN => n2302);
   U1336 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n212, B1 => 
                           REGISTERS_3_8_port, B2 => n199, ZN => n2301);
   U1337 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n238, B1 => 
                           REGISTERS_6_8_port, B2 => n225, ZN => n2300);
   U1338 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n264, B1 => 
                           REGISTERS_2_8_port, B2 => n251, ZN => n2299);
   U1339 : NAND4_X1 port map( A1 => n2302, A2 => n2301, A3 => n2300, A4 => 
                           n2299, ZN => n2308);
   U1340 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n186, B1 => 
                           REGISTERS_15_8_port, B2 => n173, ZN => n2306);
   U1341 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n212, B1 => 
                           REGISTERS_11_8_port, B2 => n199, ZN => n2305);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n238, B1 => 
                           REGISTERS_14_8_port, B2 => n225, ZN => n2304);
   U1343 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n264, B1 => 
                           REGISTERS_10_8_port, B2 => n251, ZN => n2303);
   U1344 : NAND4_X1 port map( A1 => n2306, A2 => n2305, A3 => n2304, A4 => 
                           n2303, ZN => n2307);
   U1345 : AOI22_X1 port map( A1 => n2308, A2 => n2801, B1 => n2307, B2 => 
                           n2799, ZN => n2309);
   U1346 : OAI221_X1 port map( B1 => n2805, B2 => n2311, C1 => n2803, C2 => 
                           n2310, A => n2309, ZN => N119);
   U1347 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n187, B1 => 
                           REGISTERS_23_9_port, B2 => n174, ZN => n2315);
   U1348 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n213, B1 => 
                           REGISTERS_19_9_port, B2 => n200, ZN => n2314);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n239, B1 => 
                           REGISTERS_22_9_port, B2 => n226, ZN => n2313);
   U1350 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n265, B1 => 
                           REGISTERS_18_9_port, B2 => n252, ZN => n2312);
   U1351 : AND4_X1 port map( A1 => n2315, A2 => n2314, A3 => n2313, A4 => n2312
                           , ZN => n2332);
   U1352 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n187, B1 => 
                           REGISTERS_31_9_port, B2 => n174, ZN => n2319);
   U1353 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n213, B1 => 
                           REGISTERS_27_9_port, B2 => n200, ZN => n2318);
   U1354 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n239, B1 => 
                           REGISTERS_30_9_port, B2 => n226, ZN => n2317);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n265, B1 => 
                           REGISTERS_26_9_port, B2 => n252, ZN => n2316);
   U1356 : AND4_X1 port map( A1 => n2319, A2 => n2318, A3 => n2317, A4 => n2316
                           , ZN => n2331);
   U1357 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n187, B1 => 
                           REGISTERS_7_9_port, B2 => n174, ZN => n2323);
   U1358 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n213, B1 => 
                           REGISTERS_3_9_port, B2 => n200, ZN => n2322);
   U1359 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n239, B1 => 
                           REGISTERS_6_9_port, B2 => n226, ZN => n2321);
   U1360 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n265, B1 => 
                           REGISTERS_2_9_port, B2 => n252, ZN => n2320);
   U1361 : NAND4_X1 port map( A1 => n2323, A2 => n2322, A3 => n2321, A4 => 
                           n2320, ZN => n2329);
   U1362 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n187, B1 => 
                           REGISTERS_15_9_port, B2 => n174, ZN => n2327);
   U1363 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n213, B1 => 
                           REGISTERS_11_9_port, B2 => n200, ZN => n2326);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n239, B1 => 
                           REGISTERS_14_9_port, B2 => n226, ZN => n2325);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n265, B1 => 
                           REGISTERS_10_9_port, B2 => n252, ZN => n2324);
   U1366 : NAND4_X1 port map( A1 => n2327, A2 => n2326, A3 => n2325, A4 => 
                           n2324, ZN => n2328);
   U1367 : AOI22_X1 port map( A1 => n2329, A2 => n2801, B1 => n2328, B2 => 
                           n2799, ZN => n2330);
   U1368 : OAI221_X1 port map( B1 => n2805, B2 => n2332, C1 => n2803, C2 => 
                           n2331, A => n2330, ZN => N118);
   U1369 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n187, B1 => 
                           REGISTERS_23_10_port, B2 => n174, ZN => n2336);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n213, B1 => 
                           REGISTERS_19_10_port, B2 => n200, ZN => n2335);
   U1371 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n239, B1 => 
                           REGISTERS_22_10_port, B2 => n226, ZN => n2334);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n265, B1 => 
                           REGISTERS_18_10_port, B2 => n252, ZN => n2333);
   U1373 : AND4_X1 port map( A1 => n2336, A2 => n2335, A3 => n2334, A4 => n2333
                           , ZN => n2353);
   U1374 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n187, B1 => 
                           REGISTERS_31_10_port, B2 => n174, ZN => n2340);
   U1375 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n213, B1 => 
                           REGISTERS_27_10_port, B2 => n200, ZN => n2339);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n239, B1 => 
                           REGISTERS_30_10_port, B2 => n226, ZN => n2338);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n265, B1 => 
                           REGISTERS_26_10_port, B2 => n252, ZN => n2337);
   U1378 : AND4_X1 port map( A1 => n2340, A2 => n2339, A3 => n2338, A4 => n2337
                           , ZN => n2352);
   U1379 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n187, B1 => 
                           REGISTERS_7_10_port, B2 => n174, ZN => n2344);
   U1380 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n213, B1 => 
                           REGISTERS_3_10_port, B2 => n200, ZN => n2343);
   U1381 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n239, B1 => 
                           REGISTERS_6_10_port, B2 => n226, ZN => n2342);
   U1382 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n265, B1 => 
                           REGISTERS_2_10_port, B2 => n252, ZN => n2341);
   U1383 : NAND4_X1 port map( A1 => n2344, A2 => n2343, A3 => n2342, A4 => 
                           n2341, ZN => n2350);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n187, B1 => 
                           REGISTERS_15_10_port, B2 => n174, ZN => n2348);
   U1385 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n213, B1 => 
                           REGISTERS_11_10_port, B2 => n200, ZN => n2347);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n239, B1 => 
                           REGISTERS_14_10_port, B2 => n226, ZN => n2346);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n265, B1 => 
                           REGISTERS_10_10_port, B2 => n252, ZN => n2345);
   U1388 : NAND4_X1 port map( A1 => n2348, A2 => n2347, A3 => n2346, A4 => 
                           n2345, ZN => n2349);
   U1389 : AOI22_X1 port map( A1 => n2350, A2 => n2801, B1 => n2349, B2 => 
                           n2799, ZN => n2351);
   U1390 : OAI221_X1 port map( B1 => n2805, B2 => n2353, C1 => n2803, C2 => 
                           n2352, A => n2351, ZN => N117);
   U1391 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n187, B1 => 
                           REGISTERS_23_11_port, B2 => n174, ZN => n2357);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n213, B1 => 
                           REGISTERS_19_11_port, B2 => n200, ZN => n2356);
   U1393 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n239, B1 => 
                           REGISTERS_22_11_port, B2 => n226, ZN => n2355);
   U1394 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n265, B1 => 
                           REGISTERS_18_11_port, B2 => n252, ZN => n2354);
   U1395 : AND4_X1 port map( A1 => n2357, A2 => n2356, A3 => n2355, A4 => n2354
                           , ZN => n2374);
   U1396 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n187, B1 => 
                           REGISTERS_31_11_port, B2 => n174, ZN => n2361);
   U1397 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n213, B1 => 
                           REGISTERS_27_11_port, B2 => n200, ZN => n2360);
   U1398 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n239, B1 => 
                           REGISTERS_30_11_port, B2 => n226, ZN => n2359);
   U1399 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n265, B1 => 
                           REGISTERS_26_11_port, B2 => n252, ZN => n2358);
   U1400 : AND4_X1 port map( A1 => n2361, A2 => n2360, A3 => n2359, A4 => n2358
                           , ZN => n2373);
   U1401 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n187, B1 => 
                           REGISTERS_7_11_port, B2 => n174, ZN => n2365);
   U1402 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n213, B1 => 
                           REGISTERS_3_11_port, B2 => n200, ZN => n2364);
   U1403 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n239, B1 => 
                           REGISTERS_6_11_port, B2 => n226, ZN => n2363);
   U1404 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n265, B1 => 
                           REGISTERS_2_11_port, B2 => n252, ZN => n2362);
   U1405 : NAND4_X1 port map( A1 => n2365, A2 => n2364, A3 => n2363, A4 => 
                           n2362, ZN => n2371);
   U1406 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n187, B1 => 
                           REGISTERS_15_11_port, B2 => n174, ZN => n2369);
   U1407 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n213, B1 => 
                           REGISTERS_11_11_port, B2 => n200, ZN => n2368);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n239, B1 => 
                           REGISTERS_14_11_port, B2 => n226, ZN => n2367);
   U1409 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n265, B1 => 
                           REGISTERS_10_11_port, B2 => n252, ZN => n2366);
   U1410 : NAND4_X1 port map( A1 => n2369, A2 => n2368, A3 => n2367, A4 => 
                           n2366, ZN => n2370);
   U1411 : AOI22_X1 port map( A1 => n2371, A2 => n2801, B1 => n2370, B2 => 
                           n2799, ZN => n2372);
   U1412 : OAI221_X1 port map( B1 => n2805, B2 => n2374, C1 => n2803, C2 => 
                           n2373, A => n2372, ZN => N116);
   U1413 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n188, B1 => 
                           REGISTERS_23_12_port, B2 => n175, ZN => n2378);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n214, B1 => 
                           REGISTERS_19_12_port, B2 => n201, ZN => n2377);
   U1415 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n240, B1 => 
                           REGISTERS_22_12_port, B2 => n227, ZN => n2376);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n266, B1 => 
                           REGISTERS_18_12_port, B2 => n253, ZN => n2375);
   U1417 : AND4_X1 port map( A1 => n2378, A2 => n2377, A3 => n2376, A4 => n2375
                           , ZN => n2395);
   U1418 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n188, B1 => 
                           REGISTERS_31_12_port, B2 => n175, ZN => n2382);
   U1419 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n214, B1 => 
                           REGISTERS_27_12_port, B2 => n201, ZN => n2381);
   U1420 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n240, B1 => 
                           REGISTERS_30_12_port, B2 => n227, ZN => n2380);
   U1421 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n266, B1 => 
                           REGISTERS_26_12_port, B2 => n253, ZN => n2379);
   U1422 : AND4_X1 port map( A1 => n2382, A2 => n2381, A3 => n2380, A4 => n2379
                           , ZN => n2394);
   U1423 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n188, B1 => 
                           REGISTERS_7_12_port, B2 => n175, ZN => n2386);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n214, B1 => 
                           REGISTERS_3_12_port, B2 => n201, ZN => n2385);
   U1425 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n240, B1 => 
                           REGISTERS_6_12_port, B2 => n227, ZN => n2384);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n266, B1 => 
                           REGISTERS_2_12_port, B2 => n253, ZN => n2383);
   U1427 : NAND4_X1 port map( A1 => n2386, A2 => n2385, A3 => n2384, A4 => 
                           n2383, ZN => n2392);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n188, B1 => 
                           REGISTERS_15_12_port, B2 => n175, ZN => n2390);
   U1429 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n214, B1 => 
                           REGISTERS_11_12_port, B2 => n201, ZN => n2389);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n240, B1 => 
                           REGISTERS_14_12_port, B2 => n227, ZN => n2388);
   U1431 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n266, B1 => 
                           REGISTERS_10_12_port, B2 => n253, ZN => n2387);
   U1432 : NAND4_X1 port map( A1 => n2390, A2 => n2389, A3 => n2388, A4 => 
                           n2387, ZN => n2391);
   U1433 : AOI22_X1 port map( A1 => n2392, A2 => n2801, B1 => n2391, B2 => 
                           n2799, ZN => n2393);
   U1434 : OAI221_X1 port map( B1 => n2805, B2 => n2395, C1 => n2803, C2 => 
                           n2394, A => n2393, ZN => N115);
   U1435 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n188, B1 => 
                           REGISTERS_23_13_port, B2 => n175, ZN => n2399);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n214, B1 => 
                           REGISTERS_19_13_port, B2 => n201, ZN => n2398);
   U1437 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n240, B1 => 
                           REGISTERS_22_13_port, B2 => n227, ZN => n2397);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n266, B1 => 
                           REGISTERS_18_13_port, B2 => n253, ZN => n2396);
   U1439 : AND4_X1 port map( A1 => n2399, A2 => n2398, A3 => n2397, A4 => n2396
                           , ZN => n2416);
   U1440 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n188, B1 => 
                           REGISTERS_31_13_port, B2 => n175, ZN => n2403);
   U1441 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n214, B1 => 
                           REGISTERS_27_13_port, B2 => n201, ZN => n2402);
   U1442 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n240, B1 => 
                           REGISTERS_30_13_port, B2 => n227, ZN => n2401);
   U1443 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n266, B1 => 
                           REGISTERS_26_13_port, B2 => n253, ZN => n2400);
   U1444 : AND4_X1 port map( A1 => n2403, A2 => n2402, A3 => n2401, A4 => n2400
                           , ZN => n2415);
   U1445 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n188, B1 => 
                           REGISTERS_7_13_port, B2 => n175, ZN => n2407);
   U1446 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n214, B1 => 
                           REGISTERS_3_13_port, B2 => n201, ZN => n2406);
   U1447 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n240, B1 => 
                           REGISTERS_6_13_port, B2 => n227, ZN => n2405);
   U1448 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n266, B1 => 
                           REGISTERS_2_13_port, B2 => n253, ZN => n2404);
   U1449 : NAND4_X1 port map( A1 => n2407, A2 => n2406, A3 => n2405, A4 => 
                           n2404, ZN => n2413);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n188, B1 => 
                           REGISTERS_15_13_port, B2 => n175, ZN => n2411);
   U1451 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n214, B1 => 
                           REGISTERS_11_13_port, B2 => n201, ZN => n2410);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n240, B1 => 
                           REGISTERS_14_13_port, B2 => n227, ZN => n2409);
   U1453 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n266, B1 => 
                           REGISTERS_10_13_port, B2 => n253, ZN => n2408);
   U1454 : NAND4_X1 port map( A1 => n2411, A2 => n2410, A3 => n2409, A4 => 
                           n2408, ZN => n2412);
   U1455 : AOI22_X1 port map( A1 => n2413, A2 => n2801, B1 => n2412, B2 => 
                           n2799, ZN => n2414);
   U1456 : OAI221_X1 port map( B1 => n2805, B2 => n2416, C1 => n2803, C2 => 
                           n2415, A => n2414, ZN => N114);
   U1457 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n188, B1 => 
                           REGISTERS_23_14_port, B2 => n175, ZN => n2420);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n214, B1 => 
                           REGISTERS_19_14_port, B2 => n201, ZN => n2419);
   U1459 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n240, B1 => 
                           REGISTERS_22_14_port, B2 => n227, ZN => n2418);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n266, B1 => 
                           REGISTERS_18_14_port, B2 => n253, ZN => n2417);
   U1461 : AND4_X1 port map( A1 => n2420, A2 => n2419, A3 => n2418, A4 => n2417
                           , ZN => n2437);
   U1462 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n188, B1 => 
                           REGISTERS_31_14_port, B2 => n175, ZN => n2424);
   U1463 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n214, B1 => 
                           REGISTERS_27_14_port, B2 => n201, ZN => n2423);
   U1464 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n240, B1 => 
                           REGISTERS_30_14_port, B2 => n227, ZN => n2422);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n266, B1 => 
                           REGISTERS_26_14_port, B2 => n253, ZN => n2421);
   U1466 : AND4_X1 port map( A1 => n2424, A2 => n2423, A3 => n2422, A4 => n2421
                           , ZN => n2436);
   U1467 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n188, B1 => 
                           REGISTERS_7_14_port, B2 => n175, ZN => n2428);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n214, B1 => 
                           REGISTERS_3_14_port, B2 => n201, ZN => n2427);
   U1469 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n240, B1 => 
                           REGISTERS_6_14_port, B2 => n227, ZN => n2426);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n266, B1 => 
                           REGISTERS_2_14_port, B2 => n253, ZN => n2425);
   U1471 : NAND4_X1 port map( A1 => n2428, A2 => n2427, A3 => n2426, A4 => 
                           n2425, ZN => n2434);
   U1472 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n188, B1 => 
                           REGISTERS_15_14_port, B2 => n175, ZN => n2432);
   U1473 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n214, B1 => 
                           REGISTERS_11_14_port, B2 => n201, ZN => n2431);
   U1474 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n240, B1 => 
                           REGISTERS_14_14_port, B2 => n227, ZN => n2430);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n266, B1 => 
                           REGISTERS_10_14_port, B2 => n253, ZN => n2429);
   U1476 : NAND4_X1 port map( A1 => n2432, A2 => n2431, A3 => n2430, A4 => 
                           n2429, ZN => n2433);
   U1477 : AOI22_X1 port map( A1 => n2434, A2 => n2801, B1 => n2433, B2 => 
                           n2799, ZN => n2435);
   U1478 : OAI221_X1 port map( B1 => n2805, B2 => n2437, C1 => n2803, C2 => 
                           n2436, A => n2435, ZN => N113);
   U1479 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n189, B1 => 
                           REGISTERS_23_15_port, B2 => n176, ZN => n2441);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n215, B1 => 
                           REGISTERS_19_15_port, B2 => n202, ZN => n2440);
   U1481 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n241, B1 => 
                           REGISTERS_22_15_port, B2 => n228, ZN => n2439);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n267, B1 => 
                           REGISTERS_18_15_port, B2 => n254, ZN => n2438);
   U1483 : AND4_X1 port map( A1 => n2441, A2 => n2440, A3 => n2439, A4 => n2438
                           , ZN => n2458);
   U1484 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n189, B1 => 
                           REGISTERS_31_15_port, B2 => n176, ZN => n2445);
   U1485 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n215, B1 => 
                           REGISTERS_27_15_port, B2 => n202, ZN => n2444);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n241, B1 => 
                           REGISTERS_30_15_port, B2 => n228, ZN => n2443);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n267, B1 => 
                           REGISTERS_26_15_port, B2 => n254, ZN => n2442);
   U1488 : AND4_X1 port map( A1 => n2445, A2 => n2444, A3 => n2443, A4 => n2442
                           , ZN => n2457);
   U1489 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n189, B1 => 
                           REGISTERS_7_15_port, B2 => n176, ZN => n2449);
   U1490 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n215, B1 => 
                           REGISTERS_3_15_port, B2 => n202, ZN => n2448);
   U1491 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n241, B1 => 
                           REGISTERS_6_15_port, B2 => n228, ZN => n2447);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n267, B1 => 
                           REGISTERS_2_15_port, B2 => n254, ZN => n2446);
   U1493 : NAND4_X1 port map( A1 => n2449, A2 => n2448, A3 => n2447, A4 => 
                           n2446, ZN => n2455);
   U1494 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n189, B1 => 
                           REGISTERS_15_15_port, B2 => n176, ZN => n2453);
   U1495 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n215, B1 => 
                           REGISTERS_11_15_port, B2 => n202, ZN => n2452);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n241, B1 => 
                           REGISTERS_14_15_port, B2 => n228, ZN => n2451);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n267, B1 => 
                           REGISTERS_10_15_port, B2 => n254, ZN => n2450);
   U1498 : NAND4_X1 port map( A1 => n2453, A2 => n2452, A3 => n2451, A4 => 
                           n2450, ZN => n2454);
   U1499 : AOI22_X1 port map( A1 => n2455, A2 => n2801, B1 => n2454, B2 => 
                           n2799, ZN => n2456);
   U1500 : OAI221_X1 port map( B1 => n2805, B2 => n2458, C1 => n2803, C2 => 
                           n2457, A => n2456, ZN => N112);
   U1501 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n189, B1 => 
                           REGISTERS_23_16_port, B2 => n176, ZN => n2462);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n215, B1 => 
                           REGISTERS_19_16_port, B2 => n202, ZN => n2461);
   U1503 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n241, B1 => 
                           REGISTERS_22_16_port, B2 => n228, ZN => n2460);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n267, B1 => 
                           REGISTERS_18_16_port, B2 => n254, ZN => n2459);
   U1505 : AND4_X1 port map( A1 => n2462, A2 => n2461, A3 => n2460, A4 => n2459
                           , ZN => n2479);
   U1506 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n189, B1 => 
                           REGISTERS_31_16_port, B2 => n176, ZN => n2466);
   U1507 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n215, B1 => 
                           REGISTERS_27_16_port, B2 => n202, ZN => n2465);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n241, B1 => 
                           REGISTERS_30_16_port, B2 => n228, ZN => n2464);
   U1509 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n267, B1 => 
                           REGISTERS_26_16_port, B2 => n254, ZN => n2463);
   U1510 : AND4_X1 port map( A1 => n2466, A2 => n2465, A3 => n2464, A4 => n2463
                           , ZN => n2478);
   U1511 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n189, B1 => 
                           REGISTERS_7_16_port, B2 => n176, ZN => n2470);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n215, B1 => 
                           REGISTERS_3_16_port, B2 => n202, ZN => n2469);
   U1513 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n241, B1 => 
                           REGISTERS_6_16_port, B2 => n228, ZN => n2468);
   U1514 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n267, B1 => 
                           REGISTERS_2_16_port, B2 => n254, ZN => n2467);
   U1515 : NAND4_X1 port map( A1 => n2470, A2 => n2469, A3 => n2468, A4 => 
                           n2467, ZN => n2476);
   U1516 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n189, B1 => 
                           REGISTERS_15_16_port, B2 => n176, ZN => n2474);
   U1517 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n215, B1 => 
                           REGISTERS_11_16_port, B2 => n202, ZN => n2473);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n241, B1 => 
                           REGISTERS_14_16_port, B2 => n228, ZN => n2472);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n267, B1 => 
                           REGISTERS_10_16_port, B2 => n254, ZN => n2471);
   U1520 : NAND4_X1 port map( A1 => n2474, A2 => n2473, A3 => n2472, A4 => 
                           n2471, ZN => n2475);
   U1521 : AOI22_X1 port map( A1 => n2476, A2 => n2801, B1 => n2475, B2 => 
                           n2799, ZN => n2477);
   U1522 : OAI221_X1 port map( B1 => n2805, B2 => n2479, C1 => n2803, C2 => 
                           n2478, A => n2477, ZN => N111);
   U1523 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n189, B1 => 
                           REGISTERS_23_17_port, B2 => n176, ZN => n2483);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n215, B1 => 
                           REGISTERS_19_17_port, B2 => n202, ZN => n2482);
   U1525 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n241, B1 => 
                           REGISTERS_22_17_port, B2 => n228, ZN => n2481);
   U1526 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n267, B1 => 
                           REGISTERS_18_17_port, B2 => n254, ZN => n2480);
   U1527 : AND4_X1 port map( A1 => n2483, A2 => n2482, A3 => n2481, A4 => n2480
                           , ZN => n2500);
   U1528 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n189, B1 => 
                           REGISTERS_31_17_port, B2 => n176, ZN => n2487);
   U1529 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n215, B1 => 
                           REGISTERS_27_17_port, B2 => n202, ZN => n2486);
   U1530 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n241, B1 => 
                           REGISTERS_30_17_port, B2 => n228, ZN => n2485);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n267, B1 => 
                           REGISTERS_26_17_port, B2 => n254, ZN => n2484);
   U1532 : AND4_X1 port map( A1 => n2487, A2 => n2486, A3 => n2485, A4 => n2484
                           , ZN => n2499);
   U1533 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n189, B1 => 
                           REGISTERS_7_17_port, B2 => n176, ZN => n2491);
   U1534 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n215, B1 => 
                           REGISTERS_3_17_port, B2 => n202, ZN => n2490);
   U1535 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n241, B1 => 
                           REGISTERS_6_17_port, B2 => n228, ZN => n2489);
   U1536 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n267, B1 => 
                           REGISTERS_2_17_port, B2 => n254, ZN => n2488);
   U1537 : NAND4_X1 port map( A1 => n2491, A2 => n2490, A3 => n2489, A4 => 
                           n2488, ZN => n2497);
   U1538 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n189, B1 => 
                           REGISTERS_15_17_port, B2 => n176, ZN => n2495);
   U1539 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n215, B1 => 
                           REGISTERS_11_17_port, B2 => n202, ZN => n2494);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n241, B1 => 
                           REGISTERS_14_17_port, B2 => n228, ZN => n2493);
   U1541 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n267, B1 => 
                           REGISTERS_10_17_port, B2 => n254, ZN => n2492);
   U1542 : NAND4_X1 port map( A1 => n2495, A2 => n2494, A3 => n2493, A4 => 
                           n2492, ZN => n2496);
   U1543 : AOI22_X1 port map( A1 => n2497, A2 => n2801, B1 => n2496, B2 => 
                           n2799, ZN => n2498);
   U1544 : OAI221_X1 port map( B1 => n2805, B2 => n2500, C1 => n2803, C2 => 
                           n2499, A => n2498, ZN => N110);
   U1545 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n190, B1 => 
                           REGISTERS_23_18_port, B2 => n177, ZN => n2504);
   U1546 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n216, B1 => 
                           REGISTERS_19_18_port, B2 => n203, ZN => n2503);
   U1547 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n242, B1 => 
                           REGISTERS_22_18_port, B2 => n229, ZN => n2502);
   U1548 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n268, B1 => 
                           REGISTERS_18_18_port, B2 => n255, ZN => n2501);
   U1549 : AND4_X1 port map( A1 => n2504, A2 => n2503, A3 => n2502, A4 => n2501
                           , ZN => n2521);
   U1550 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n190, B1 => 
                           REGISTERS_31_18_port, B2 => n177, ZN => n2508);
   U1551 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n216, B1 => 
                           REGISTERS_27_18_port, B2 => n203, ZN => n2507);
   U1552 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n242, B1 => 
                           REGISTERS_30_18_port, B2 => n229, ZN => n2506);
   U1553 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n268, B1 => 
                           REGISTERS_26_18_port, B2 => n255, ZN => n2505);
   U1554 : AND4_X1 port map( A1 => n2508, A2 => n2507, A3 => n2506, A4 => n2505
                           , ZN => n2520);
   U1555 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n190, B1 => 
                           REGISTERS_7_18_port, B2 => n177, ZN => n2512);
   U1556 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n216, B1 => 
                           REGISTERS_3_18_port, B2 => n203, ZN => n2511);
   U1557 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n242, B1 => 
                           REGISTERS_6_18_port, B2 => n229, ZN => n2510);
   U1558 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n268, B1 => 
                           REGISTERS_2_18_port, B2 => n255, ZN => n2509);
   U1559 : NAND4_X1 port map( A1 => n2512, A2 => n2511, A3 => n2510, A4 => 
                           n2509, ZN => n2518);
   U1560 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n190, B1 => 
                           REGISTERS_15_18_port, B2 => n177, ZN => n2516);
   U1561 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n216, B1 => 
                           REGISTERS_11_18_port, B2 => n203, ZN => n2515);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n242, B1 => 
                           REGISTERS_14_18_port, B2 => n229, ZN => n2514);
   U1563 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n268, B1 => 
                           REGISTERS_10_18_port, B2 => n255, ZN => n2513);
   U1564 : NAND4_X1 port map( A1 => n2516, A2 => n2515, A3 => n2514, A4 => 
                           n2513, ZN => n2517);
   U1565 : AOI22_X1 port map( A1 => n2518, A2 => n2801, B1 => n2517, B2 => 
                           n2799, ZN => n2519);
   U1566 : OAI221_X1 port map( B1 => n2805, B2 => n2521, C1 => n2803, C2 => 
                           n2520, A => n2519, ZN => N109);
   U1567 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n190, B1 => 
                           REGISTERS_23_19_port, B2 => n177, ZN => n2525);
   U1568 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n216, B1 => 
                           REGISTERS_19_19_port, B2 => n203, ZN => n2524);
   U1569 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n242, B1 => 
                           REGISTERS_22_19_port, B2 => n229, ZN => n2523);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n268, B1 => 
                           REGISTERS_18_19_port, B2 => n255, ZN => n2522);
   U1571 : AND4_X1 port map( A1 => n2525, A2 => n2524, A3 => n2523, A4 => n2522
                           , ZN => n2542);
   U1572 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n190, B1 => 
                           REGISTERS_31_19_port, B2 => n177, ZN => n2529);
   U1573 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n216, B1 => 
                           REGISTERS_27_19_port, B2 => n203, ZN => n2528);
   U1574 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n242, B1 => 
                           REGISTERS_30_19_port, B2 => n229, ZN => n2527);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n268, B1 => 
                           REGISTERS_26_19_port, B2 => n255, ZN => n2526);
   U1576 : AND4_X1 port map( A1 => n2529, A2 => n2528, A3 => n2527, A4 => n2526
                           , ZN => n2541);
   U1577 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n190, B1 => 
                           REGISTERS_7_19_port, B2 => n177, ZN => n2533);
   U1578 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n216, B1 => 
                           REGISTERS_3_19_port, B2 => n203, ZN => n2532);
   U1579 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n242, B1 => 
                           REGISTERS_6_19_port, B2 => n229, ZN => n2531);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n268, B1 => 
                           REGISTERS_2_19_port, B2 => n255, ZN => n2530);
   U1581 : NAND4_X1 port map( A1 => n2533, A2 => n2532, A3 => n2531, A4 => 
                           n2530, ZN => n2539);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n190, B1 => 
                           REGISTERS_15_19_port, B2 => n177, ZN => n2537);
   U1583 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n216, B1 => 
                           REGISTERS_11_19_port, B2 => n203, ZN => n2536);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n242, B1 => 
                           REGISTERS_14_19_port, B2 => n229, ZN => n2535);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n268, B1 => 
                           REGISTERS_10_19_port, B2 => n255, ZN => n2534);
   U1586 : NAND4_X1 port map( A1 => n2537, A2 => n2536, A3 => n2535, A4 => 
                           n2534, ZN => n2538);
   U1587 : AOI22_X1 port map( A1 => n2539, A2 => n2801, B1 => n2538, B2 => 
                           n2799, ZN => n2540);
   U1588 : OAI221_X1 port map( B1 => n2805, B2 => n2542, C1 => n2803, C2 => 
                           n2541, A => n2540, ZN => N108);
   U1589 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n190, B1 => 
                           REGISTERS_23_20_port, B2 => n177, ZN => n2546);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n216, B1 => 
                           REGISTERS_19_20_port, B2 => n203, ZN => n2545);
   U1591 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n242, B1 => 
                           REGISTERS_22_20_port, B2 => n229, ZN => n2544);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n268, B1 => 
                           REGISTERS_18_20_port, B2 => n255, ZN => n2543);
   U1593 : AND4_X1 port map( A1 => n2546, A2 => n2545, A3 => n2544, A4 => n2543
                           , ZN => n2563);
   U1594 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n190, B1 => 
                           REGISTERS_31_20_port, B2 => n177, ZN => n2550);
   U1595 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n216, B1 => 
                           REGISTERS_27_20_port, B2 => n203, ZN => n2549);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n242, B1 => 
                           REGISTERS_30_20_port, B2 => n229, ZN => n2548);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n268, B1 => 
                           REGISTERS_26_20_port, B2 => n255, ZN => n2547);
   U1598 : AND4_X1 port map( A1 => n2550, A2 => n2549, A3 => n2548, A4 => n2547
                           , ZN => n2562);
   U1599 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n190, B1 => 
                           REGISTERS_7_20_port, B2 => n177, ZN => n2554);
   U1600 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n216, B1 => 
                           REGISTERS_3_20_port, B2 => n203, ZN => n2553);
   U1601 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n242, B1 => 
                           REGISTERS_6_20_port, B2 => n229, ZN => n2552);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n268, B1 => 
                           REGISTERS_2_20_port, B2 => n255, ZN => n2551);
   U1603 : NAND4_X1 port map( A1 => n2554, A2 => n2553, A3 => n2552, A4 => 
                           n2551, ZN => n2560);
   U1604 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n190, B1 => 
                           REGISTERS_15_20_port, B2 => n177, ZN => n2558);
   U1605 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n216, B1 => 
                           REGISTERS_11_20_port, B2 => n203, ZN => n2557);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n242, B1 => 
                           REGISTERS_14_20_port, B2 => n229, ZN => n2556);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n268, B1 => 
                           REGISTERS_10_20_port, B2 => n255, ZN => n2555);
   U1608 : NAND4_X1 port map( A1 => n2558, A2 => n2557, A3 => n2556, A4 => 
                           n2555, ZN => n2559);
   U1609 : AOI22_X1 port map( A1 => n2560, A2 => n2801, B1 => n2559, B2 => 
                           n2799, ZN => n2561);
   U1610 : OAI221_X1 port map( B1 => n2805, B2 => n2563, C1 => n2803, C2 => 
                           n2562, A => n2561, ZN => N107);
   U1611 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n191, B1 => 
                           REGISTERS_23_21_port, B2 => n178, ZN => n2567);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n217, B1 => 
                           REGISTERS_19_21_port, B2 => n204, ZN => n2566);
   U1613 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n243, B1 => 
                           REGISTERS_22_21_port, B2 => n230, ZN => n2565);
   U1614 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n269, B1 => 
                           REGISTERS_18_21_port, B2 => n256, ZN => n2564);
   U1615 : AND4_X1 port map( A1 => n2567, A2 => n2566, A3 => n2565, A4 => n2564
                           , ZN => n2584);
   U1616 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n191, B1 => 
                           REGISTERS_31_21_port, B2 => n178, ZN => n2571);
   U1617 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n217, B1 => 
                           REGISTERS_27_21_port, B2 => n204, ZN => n2570);
   U1618 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n243, B1 => 
                           REGISTERS_30_21_port, B2 => n230, ZN => n2569);
   U1619 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n269, B1 => 
                           REGISTERS_26_21_port, B2 => n256, ZN => n2568);
   U1620 : AND4_X1 port map( A1 => n2571, A2 => n2570, A3 => n2569, A4 => n2568
                           , ZN => n2583);
   U1621 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n191, B1 => 
                           REGISTERS_7_21_port, B2 => n178, ZN => n2575);
   U1622 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n217, B1 => 
                           REGISTERS_3_21_port, B2 => n204, ZN => n2574);
   U1623 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n243, B1 => 
                           REGISTERS_6_21_port, B2 => n230, ZN => n2573);
   U1624 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n269, B1 => 
                           REGISTERS_2_21_port, B2 => n256, ZN => n2572);
   U1625 : NAND4_X1 port map( A1 => n2575, A2 => n2574, A3 => n2573, A4 => 
                           n2572, ZN => n2581);
   U1626 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n191, B1 => 
                           REGISTERS_15_21_port, B2 => n178, ZN => n2579);
   U1627 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n217, B1 => 
                           REGISTERS_11_21_port, B2 => n204, ZN => n2578);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n243, B1 => 
                           REGISTERS_14_21_port, B2 => n230, ZN => n2577);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n269, B1 => 
                           REGISTERS_10_21_port, B2 => n256, ZN => n2576);
   U1630 : NAND4_X1 port map( A1 => n2579, A2 => n2578, A3 => n2577, A4 => 
                           n2576, ZN => n2580);
   U1631 : AOI22_X1 port map( A1 => n2581, A2 => n2801, B1 => n2580, B2 => 
                           n2799, ZN => n2582);
   U1632 : OAI221_X1 port map( B1 => n2805, B2 => n2584, C1 => n2803, C2 => 
                           n2583, A => n2582, ZN => N106);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n191, B1 => 
                           REGISTERS_23_22_port, B2 => n178, ZN => n2588);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n217, B1 => 
                           REGISTERS_19_22_port, B2 => n204, ZN => n2587);
   U1635 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n243, B1 => 
                           REGISTERS_22_22_port, B2 => n230, ZN => n2586);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n269, B1 => 
                           REGISTERS_18_22_port, B2 => n256, ZN => n2585);
   U1637 : AND4_X1 port map( A1 => n2588, A2 => n2587, A3 => n2586, A4 => n2585
                           , ZN => n2605);
   U1638 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n191, B1 => 
                           REGISTERS_31_22_port, B2 => n178, ZN => n2592);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n217, B1 => 
                           REGISTERS_27_22_port, B2 => n204, ZN => n2591);
   U1640 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n243, B1 => 
                           REGISTERS_30_22_port, B2 => n230, ZN => n2590);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n269, B1 => 
                           REGISTERS_26_22_port, B2 => n256, ZN => n2589);
   U1642 : AND4_X1 port map( A1 => n2592, A2 => n2591, A3 => n2590, A4 => n2589
                           , ZN => n2604);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n191, B1 => 
                           REGISTERS_7_22_port, B2 => n178, ZN => n2596);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n217, B1 => 
                           REGISTERS_3_22_port, B2 => n204, ZN => n2595);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n243, B1 => 
                           REGISTERS_6_22_port, B2 => n230, ZN => n2594);
   U1646 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n269, B1 => 
                           REGISTERS_2_22_port, B2 => n256, ZN => n2593);
   U1647 : NAND4_X1 port map( A1 => n2596, A2 => n2595, A3 => n2594, A4 => 
                           n2593, ZN => n2602);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n191, B1 => 
                           REGISTERS_15_22_port, B2 => n178, ZN => n2600);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n217, B1 => 
                           REGISTERS_11_22_port, B2 => n204, ZN => n2599);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n243, B1 => 
                           REGISTERS_14_22_port, B2 => n230, ZN => n2598);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n269, B1 => 
                           REGISTERS_10_22_port, B2 => n256, ZN => n2597);
   U1652 : NAND4_X1 port map( A1 => n2600, A2 => n2599, A3 => n2598, A4 => 
                           n2597, ZN => n2601);
   U1653 : AOI22_X1 port map( A1 => n2602, A2 => n2801, B1 => n2601, B2 => 
                           n2799, ZN => n2603);
   U1654 : OAI221_X1 port map( B1 => n2805, B2 => n2605, C1 => n2803, C2 => 
                           n2604, A => n2603, ZN => N105);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n191, B1 => 
                           REGISTERS_23_23_port, B2 => n178, ZN => n2609);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n217, B1 => 
                           REGISTERS_19_23_port, B2 => n204, ZN => n2608);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n243, B1 => 
                           REGISTERS_22_23_port, B2 => n230, ZN => n2607);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n269, B1 => 
                           REGISTERS_18_23_port, B2 => n256, ZN => n2606);
   U1659 : AND4_X1 port map( A1 => n2609, A2 => n2608, A3 => n2607, A4 => n2606
                           , ZN => n2626);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n191, B1 => 
                           REGISTERS_31_23_port, B2 => n178, ZN => n2613);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n217, B1 => 
                           REGISTERS_27_23_port, B2 => n204, ZN => n2612);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n243, B1 => 
                           REGISTERS_30_23_port, B2 => n230, ZN => n2611);
   U1663 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n269, B1 => 
                           REGISTERS_26_23_port, B2 => n256, ZN => n2610);
   U1664 : AND4_X1 port map( A1 => n2613, A2 => n2612, A3 => n2611, A4 => n2610
                           , ZN => n2625);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n191, B1 => 
                           REGISTERS_7_23_port, B2 => n178, ZN => n2617);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n217, B1 => 
                           REGISTERS_3_23_port, B2 => n204, ZN => n2616);
   U1667 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n243, B1 => 
                           REGISTERS_6_23_port, B2 => n230, ZN => n2615);
   U1668 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n269, B1 => 
                           REGISTERS_2_23_port, B2 => n256, ZN => n2614);
   U1669 : NAND4_X1 port map( A1 => n2617, A2 => n2616, A3 => n2615, A4 => 
                           n2614, ZN => n2623);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n191, B1 => 
                           REGISTERS_15_23_port, B2 => n178, ZN => n2621);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n217, B1 => 
                           REGISTERS_11_23_port, B2 => n204, ZN => n2620);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n243, B1 => 
                           REGISTERS_14_23_port, B2 => n230, ZN => n2619);
   U1673 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n269, B1 => 
                           REGISTERS_10_23_port, B2 => n256, ZN => n2618);
   U1674 : NAND4_X1 port map( A1 => n2621, A2 => n2620, A3 => n2619, A4 => 
                           n2618, ZN => n2622);
   U1675 : AOI22_X1 port map( A1 => n2623, A2 => n2801, B1 => n2622, B2 => 
                           n2799, ZN => n2624);
   U1676 : OAI221_X1 port map( B1 => n2805, B2 => n2626, C1 => n2803, C2 => 
                           n2625, A => n2624, ZN => N104);
   U1677 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n192, B1 => 
                           REGISTERS_23_24_port, B2 => n179, ZN => n2630);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n218, B1 => 
                           REGISTERS_19_24_port, B2 => n205, ZN => n2629);
   U1679 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n244, B1 => 
                           REGISTERS_22_24_port, B2 => n231, ZN => n2628);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n270, B1 => 
                           REGISTERS_18_24_port, B2 => n257, ZN => n2627);
   U1681 : AND4_X1 port map( A1 => n2630, A2 => n2629, A3 => n2628, A4 => n2627
                           , ZN => n2647);
   U1682 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n192, B1 => 
                           REGISTERS_31_24_port, B2 => n179, ZN => n2634);
   U1683 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n218, B1 => 
                           REGISTERS_27_24_port, B2 => n205, ZN => n2633);
   U1684 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n244, B1 => 
                           REGISTERS_30_24_port, B2 => n231, ZN => n2632);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n270, B1 => 
                           REGISTERS_26_24_port, B2 => n257, ZN => n2631);
   U1686 : AND4_X1 port map( A1 => n2634, A2 => n2633, A3 => n2632, A4 => n2631
                           , ZN => n2646);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n192, B1 => 
                           REGISTERS_7_24_port, B2 => n179, ZN => n2638);
   U1688 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n218, B1 => 
                           REGISTERS_3_24_port, B2 => n205, ZN => n2637);
   U1689 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n244, B1 => 
                           REGISTERS_6_24_port, B2 => n231, ZN => n2636);
   U1690 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n270, B1 => 
                           REGISTERS_2_24_port, B2 => n257, ZN => n2635);
   U1691 : NAND4_X1 port map( A1 => n2638, A2 => n2637, A3 => n2636, A4 => 
                           n2635, ZN => n2644);
   U1692 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n192, B1 => 
                           REGISTERS_15_24_port, B2 => n179, ZN => n2642);
   U1693 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n218, B1 => 
                           REGISTERS_11_24_port, B2 => n205, ZN => n2641);
   U1694 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n244, B1 => 
                           REGISTERS_14_24_port, B2 => n231, ZN => n2640);
   U1695 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n270, B1 => 
                           REGISTERS_10_24_port, B2 => n257, ZN => n2639);
   U1696 : NAND4_X1 port map( A1 => n2642, A2 => n2641, A3 => n2640, A4 => 
                           n2639, ZN => n2643);
   U1697 : AOI22_X1 port map( A1 => n2644, A2 => n2801, B1 => n2643, B2 => 
                           n2799, ZN => n2645);
   U1698 : OAI221_X1 port map( B1 => n2805, B2 => n2647, C1 => n2803, C2 => 
                           n2646, A => n2645, ZN => N103);
   U1699 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n192, B1 => 
                           REGISTERS_23_25_port, B2 => n179, ZN => n2651);
   U1700 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n218, B1 => 
                           REGISTERS_19_25_port, B2 => n205, ZN => n2650);
   U1701 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n244, B1 => 
                           REGISTERS_22_25_port, B2 => n231, ZN => n2649);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n270, B1 => 
                           REGISTERS_18_25_port, B2 => n257, ZN => n2648);
   U1703 : AND4_X1 port map( A1 => n2651, A2 => n2650, A3 => n2649, A4 => n2648
                           , ZN => n2668);
   U1704 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n192, B1 => 
                           REGISTERS_31_25_port, B2 => n179, ZN => n2655);
   U1705 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n218, B1 => 
                           REGISTERS_27_25_port, B2 => n205, ZN => n2654);
   U1706 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n244, B1 => 
                           REGISTERS_30_25_port, B2 => n231, ZN => n2653);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n270, B1 => 
                           REGISTERS_26_25_port, B2 => n257, ZN => n2652);
   U1708 : AND4_X1 port map( A1 => n2655, A2 => n2654, A3 => n2653, A4 => n2652
                           , ZN => n2667);
   U1709 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n192, B1 => 
                           REGISTERS_7_25_port, B2 => n179, ZN => n2659);
   U1710 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n218, B1 => 
                           REGISTERS_3_25_port, B2 => n205, ZN => n2658);
   U1711 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n244, B1 => 
                           REGISTERS_6_25_port, B2 => n231, ZN => n2657);
   U1712 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n270, B1 => 
                           REGISTERS_2_25_port, B2 => n257, ZN => n2656);
   U1713 : NAND4_X1 port map( A1 => n2659, A2 => n2658, A3 => n2657, A4 => 
                           n2656, ZN => n2665);
   U1714 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n192, B1 => 
                           REGISTERS_15_25_port, B2 => n179, ZN => n2663);
   U1715 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n218, B1 => 
                           REGISTERS_11_25_port, B2 => n205, ZN => n2662);
   U1716 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n244, B1 => 
                           REGISTERS_14_25_port, B2 => n231, ZN => n2661);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n270, B1 => 
                           REGISTERS_10_25_port, B2 => n257, ZN => n2660);
   U1718 : NAND4_X1 port map( A1 => n2663, A2 => n2662, A3 => n2661, A4 => 
                           n2660, ZN => n2664);
   U1719 : AOI22_X1 port map( A1 => n2665, A2 => n2801, B1 => n2664, B2 => 
                           n2799, ZN => n2666);
   U1720 : OAI221_X1 port map( B1 => n2805, B2 => n2668, C1 => n2803, C2 => 
                           n2667, A => n2666, ZN => N102);
   U1721 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n192, B1 => 
                           REGISTERS_23_26_port, B2 => n179, ZN => n2672);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n218, B1 => 
                           REGISTERS_19_26_port, B2 => n205, ZN => n2671);
   U1723 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n244, B1 => 
                           REGISTERS_22_26_port, B2 => n231, ZN => n2670);
   U1724 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n270, B1 => 
                           REGISTERS_18_26_port, B2 => n257, ZN => n2669);
   U1725 : AND4_X1 port map( A1 => n2672, A2 => n2671, A3 => n2670, A4 => n2669
                           , ZN => n2689);
   U1726 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n192, B1 => 
                           REGISTERS_31_26_port, B2 => n179, ZN => n2676);
   U1727 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n218, B1 => 
                           REGISTERS_27_26_port, B2 => n205, ZN => n2675);
   U1728 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n244, B1 => 
                           REGISTERS_30_26_port, B2 => n231, ZN => n2674);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n270, B1 => 
                           REGISTERS_26_26_port, B2 => n257, ZN => n2673);
   U1730 : AND4_X1 port map( A1 => n2676, A2 => n2675, A3 => n2674, A4 => n2673
                           , ZN => n2688);
   U1731 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n192, B1 => 
                           REGISTERS_7_26_port, B2 => n179, ZN => n2680);
   U1732 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n218, B1 => 
                           REGISTERS_3_26_port, B2 => n205, ZN => n2679);
   U1733 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n244, B1 => 
                           REGISTERS_6_26_port, B2 => n231, ZN => n2678);
   U1734 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n270, B1 => 
                           REGISTERS_2_26_port, B2 => n257, ZN => n2677);
   U1735 : NAND4_X1 port map( A1 => n2680, A2 => n2679, A3 => n2678, A4 => 
                           n2677, ZN => n2686);
   U1736 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n192, B1 => 
                           REGISTERS_15_26_port, B2 => n179, ZN => n2684);
   U1737 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n218, B1 => 
                           REGISTERS_11_26_port, B2 => n205, ZN => n2683);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n244, B1 => 
                           REGISTERS_14_26_port, B2 => n231, ZN => n2682);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n270, B1 => 
                           REGISTERS_10_26_port, B2 => n257, ZN => n2681);
   U1740 : NAND4_X1 port map( A1 => n2684, A2 => n2683, A3 => n2682, A4 => 
                           n2681, ZN => n2685);
   U1741 : AOI22_X1 port map( A1 => n2686, A2 => n2801, B1 => n2685, B2 => 
                           n2799, ZN => n2687);
   U1742 : OAI221_X1 port map( B1 => n2805, B2 => n2689, C1 => n2803, C2 => 
                           n2688, A => n2687, ZN => N101);
   U1743 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n193, B1 => 
                           REGISTERS_23_27_port, B2 => n180, ZN => n2693);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n219, B1 => 
                           REGISTERS_19_27_port, B2 => n206, ZN => n2692);
   U1745 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n245, B1 => 
                           REGISTERS_22_27_port, B2 => n232, ZN => n2691);
   U1746 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n271, B1 => 
                           REGISTERS_18_27_port, B2 => n258, ZN => n2690);
   U1747 : AND4_X1 port map( A1 => n2693, A2 => n2692, A3 => n2691, A4 => n2690
                           , ZN => n2710);
   U1748 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n193, B1 => 
                           REGISTERS_31_27_port, B2 => n180, ZN => n2697);
   U1749 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n219, B1 => 
                           REGISTERS_27_27_port, B2 => n206, ZN => n2696);
   U1750 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n245, B1 => 
                           REGISTERS_30_27_port, B2 => n232, ZN => n2695);
   U1751 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n271, B1 => 
                           REGISTERS_26_27_port, B2 => n258, ZN => n2694);
   U1752 : AND4_X1 port map( A1 => n2697, A2 => n2696, A3 => n2695, A4 => n2694
                           , ZN => n2709);
   U1753 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n193, B1 => 
                           REGISTERS_7_27_port, B2 => n180, ZN => n2701);
   U1754 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n219, B1 => 
                           REGISTERS_3_27_port, B2 => n206, ZN => n2700);
   U1755 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n245, B1 => 
                           REGISTERS_6_27_port, B2 => n232, ZN => n2699);
   U1756 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n271, B1 => 
                           REGISTERS_2_27_port, B2 => n258, ZN => n2698);
   U1757 : NAND4_X1 port map( A1 => n2701, A2 => n2700, A3 => n2699, A4 => 
                           n2698, ZN => n2707);
   U1758 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n193, B1 => 
                           REGISTERS_15_27_port, B2 => n180, ZN => n2705);
   U1759 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n219, B1 => 
                           REGISTERS_11_27_port, B2 => n206, ZN => n2704);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n245, B1 => 
                           REGISTERS_14_27_port, B2 => n232, ZN => n2703);
   U1761 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n271, B1 => 
                           REGISTERS_10_27_port, B2 => n258, ZN => n2702);
   U1762 : NAND4_X1 port map( A1 => n2705, A2 => n2704, A3 => n2703, A4 => 
                           n2702, ZN => n2706);
   U1763 : AOI22_X1 port map( A1 => n2707, A2 => n2801, B1 => n2706, B2 => 
                           n2799, ZN => n2708);
   U1764 : OAI221_X1 port map( B1 => n2805, B2 => n2710, C1 => n2803, C2 => 
                           n2709, A => n2708, ZN => N100);
   U1765 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n193, B1 => 
                           REGISTERS_23_28_port, B2 => n180, ZN => n2714);
   U1766 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n219, B1 => 
                           REGISTERS_19_28_port, B2 => n206, ZN => n2713);
   U1767 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n245, B1 => 
                           REGISTERS_22_28_port, B2 => n232, ZN => n2712);
   U1768 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n271, B1 => 
                           REGISTERS_18_28_port, B2 => n258, ZN => n2711);
   U1769 : AND4_X1 port map( A1 => n2714, A2 => n2713, A3 => n2712, A4 => n2711
                           , ZN => n2731);
   U1770 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n193, B1 => 
                           REGISTERS_31_28_port, B2 => n180, ZN => n2718);
   U1771 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n219, B1 => 
                           REGISTERS_27_28_port, B2 => n206, ZN => n2717);
   U1772 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n245, B1 => 
                           REGISTERS_30_28_port, B2 => n232, ZN => n2716);
   U1773 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n271, B1 => 
                           REGISTERS_26_28_port, B2 => n258, ZN => n2715);
   U1774 : AND4_X1 port map( A1 => n2718, A2 => n2717, A3 => n2716, A4 => n2715
                           , ZN => n2730);
   U1775 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n193, B1 => 
                           REGISTERS_7_28_port, B2 => n180, ZN => n2722);
   U1776 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n219, B1 => 
                           REGISTERS_3_28_port, B2 => n206, ZN => n2721);
   U1777 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n245, B1 => 
                           REGISTERS_6_28_port, B2 => n232, ZN => n2720);
   U1778 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n271, B1 => 
                           REGISTERS_2_28_port, B2 => n258, ZN => n2719);
   U1779 : NAND4_X1 port map( A1 => n2722, A2 => n2721, A3 => n2720, A4 => 
                           n2719, ZN => n2728);
   U1780 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n193, B1 => 
                           REGISTERS_15_28_port, B2 => n180, ZN => n2726);
   U1781 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n219, B1 => 
                           REGISTERS_11_28_port, B2 => n206, ZN => n2725);
   U1782 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n245, B1 => 
                           REGISTERS_14_28_port, B2 => n232, ZN => n2724);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n271, B1 => 
                           REGISTERS_10_28_port, B2 => n258, ZN => n2723);
   U1784 : NAND4_X1 port map( A1 => n2726, A2 => n2725, A3 => n2724, A4 => 
                           n2723, ZN => n2727);
   U1785 : AOI22_X1 port map( A1 => n2728, A2 => n2801, B1 => n2727, B2 => 
                           n2799, ZN => n2729);
   U1786 : OAI221_X1 port map( B1 => n2805, B2 => n2731, C1 => n2803, C2 => 
                           n2730, A => n2729, ZN => N99);
   U1787 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n193, B1 => 
                           REGISTERS_23_29_port, B2 => n180, ZN => n2735);
   U1788 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n219, B1 => 
                           REGISTERS_19_29_port, B2 => n206, ZN => n2734);
   U1789 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n245, B1 => 
                           REGISTERS_22_29_port, B2 => n232, ZN => n2733);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n271, B1 => 
                           REGISTERS_18_29_port, B2 => n258, ZN => n2732);
   U1791 : AND4_X1 port map( A1 => n2735, A2 => n2734, A3 => n2733, A4 => n2732
                           , ZN => n2752);
   U1792 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n193, B1 => 
                           REGISTERS_31_29_port, B2 => n180, ZN => n2739);
   U1793 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n219, B1 => 
                           REGISTERS_27_29_port, B2 => n206, ZN => n2738);
   U1794 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n245, B1 => 
                           REGISTERS_30_29_port, B2 => n232, ZN => n2737);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n271, B1 => 
                           REGISTERS_26_29_port, B2 => n258, ZN => n2736);
   U1796 : AND4_X1 port map( A1 => n2739, A2 => n2738, A3 => n2737, A4 => n2736
                           , ZN => n2751);
   U1797 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n193, B1 => 
                           REGISTERS_7_29_port, B2 => n180, ZN => n2743);
   U1798 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n219, B1 => 
                           REGISTERS_3_29_port, B2 => n206, ZN => n2742);
   U1799 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n245, B1 => 
                           REGISTERS_6_29_port, B2 => n232, ZN => n2741);
   U1800 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n271, B1 => 
                           REGISTERS_2_29_port, B2 => n258, ZN => n2740);
   U1801 : NAND4_X1 port map( A1 => n2743, A2 => n2742, A3 => n2741, A4 => 
                           n2740, ZN => n2749);
   U1802 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n193, B1 => 
                           REGISTERS_15_29_port, B2 => n180, ZN => n2747);
   U1803 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n219, B1 => 
                           REGISTERS_11_29_port, B2 => n206, ZN => n2746);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n245, B1 => 
                           REGISTERS_14_29_port, B2 => n232, ZN => n2745);
   U1805 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n271, B1 => 
                           REGISTERS_10_29_port, B2 => n258, ZN => n2744);
   U1806 : NAND4_X1 port map( A1 => n2747, A2 => n2746, A3 => n2745, A4 => 
                           n2744, ZN => n2748);
   U1807 : AOI22_X1 port map( A1 => n2749, A2 => n2801, B1 => n2748, B2 => 
                           n2799, ZN => n2750);
   U1808 : OAI221_X1 port map( B1 => n2805, B2 => n2752, C1 => n2803, C2 => 
                           n2751, A => n2750, ZN => N98);
   U1809 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n194, B1 => 
                           REGISTERS_23_30_port, B2 => n181, ZN => n2756);
   U1810 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n220, B1 => 
                           REGISTERS_19_30_port, B2 => n207, ZN => n2755);
   U1811 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n246, B1 => 
                           REGISTERS_22_30_port, B2 => n233, ZN => n2754);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n272, B1 => 
                           REGISTERS_18_30_port, B2 => n259, ZN => n2753);
   U1813 : AND4_X1 port map( A1 => n2756, A2 => n2755, A3 => n2754, A4 => n2753
                           , ZN => n2773);
   U1814 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n194, B1 => 
                           REGISTERS_31_30_port, B2 => n181, ZN => n2760);
   U1815 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n220, B1 => 
                           REGISTERS_27_30_port, B2 => n207, ZN => n2759);
   U1816 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n246, B1 => 
                           REGISTERS_30_30_port, B2 => n233, ZN => n2758);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n272, B1 => 
                           REGISTERS_26_30_port, B2 => n259, ZN => n2757);
   U1818 : AND4_X1 port map( A1 => n2760, A2 => n2759, A3 => n2758, A4 => n2757
                           , ZN => n2772);
   U1819 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n194, B1 => 
                           REGISTERS_7_30_port, B2 => n181, ZN => n2764);
   U1820 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n220, B1 => 
                           REGISTERS_3_30_port, B2 => n207, ZN => n2763);
   U1821 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n246, B1 => 
                           REGISTERS_6_30_port, B2 => n233, ZN => n2762);
   U1822 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n272, B1 => 
                           REGISTERS_2_30_port, B2 => n259, ZN => n2761);
   U1823 : NAND4_X1 port map( A1 => n2764, A2 => n2763, A3 => n2762, A4 => 
                           n2761, ZN => n2770);
   U1824 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n194, B1 => 
                           REGISTERS_15_30_port, B2 => n181, ZN => n2768);
   U1825 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n220, B1 => 
                           REGISTERS_11_30_port, B2 => n207, ZN => n2767);
   U1826 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n246, B1 => 
                           REGISTERS_14_30_port, B2 => n233, ZN => n2766);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n272, B1 => 
                           REGISTERS_10_30_port, B2 => n259, ZN => n2765);
   U1828 : NAND4_X1 port map( A1 => n2768, A2 => n2767, A3 => n2766, A4 => 
                           n2765, ZN => n2769);
   U1829 : AOI22_X1 port map( A1 => n2770, A2 => n2801, B1 => n2769, B2 => 
                           n2799, ZN => n2771);
   U1830 : OAI221_X1 port map( B1 => n2805, B2 => n2773, C1 => n2803, C2 => 
                           n2772, A => n2771, ZN => N97);
   U1831 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n194, B1 => 
                           REGISTERS_23_31_port, B2 => n181, ZN => n2777);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n220, B1 => 
                           REGISTERS_19_31_port, B2 => n207, ZN => n2776);
   U1833 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n246, B1 => 
                           REGISTERS_22_31_port, B2 => n233, ZN => n2775);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n272, B1 => 
                           REGISTERS_18_31_port, B2 => n259, ZN => n2774);
   U1835 : AND4_X1 port map( A1 => n2777, A2 => n2776, A3 => n2775, A4 => n2774
                           , ZN => n2806);
   U1836 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n194, B1 => 
                           REGISTERS_31_31_port, B2 => n181, ZN => n2781);
   U1837 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n220, B1 => 
                           REGISTERS_27_31_port, B2 => n207, ZN => n2780);
   U1838 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n246, B1 => 
                           REGISTERS_30_31_port, B2 => n233, ZN => n2779);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n272, B1 => 
                           REGISTERS_26_31_port, B2 => n259, ZN => n2778);
   U1840 : AND4_X1 port map( A1 => n2781, A2 => n2780, A3 => n2779, A4 => n2778
                           , ZN => n2804);
   U1841 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n194, B1 => 
                           REGISTERS_7_31_port, B2 => n181, ZN => n2785);
   U1842 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n220, B1 => 
                           REGISTERS_3_31_port, B2 => n207, ZN => n2784);
   U1843 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n246, B1 => 
                           REGISTERS_6_31_port, B2 => n233, ZN => n2783);
   U1844 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n272, B1 => 
                           REGISTERS_2_31_port, B2 => n259, ZN => n2782);
   U1845 : NAND4_X1 port map( A1 => n2785, A2 => n2784, A3 => n2783, A4 => 
                           n2782, ZN => n2800);
   U1846 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n194, B1 => 
                           REGISTERS_15_31_port, B2 => n181, ZN => n2797);
   U1847 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n220, B1 => 
                           REGISTERS_11_31_port, B2 => n207, ZN => n2796);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n246, B1 => 
                           REGISTERS_14_31_port, B2 => n233, ZN => n2795);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n272, B1 => 
                           REGISTERS_10_31_port, B2 => n259, ZN => n2794);
   U1850 : NAND4_X1 port map( A1 => n2797, A2 => n2796, A3 => n2795, A4 => 
                           n2794, ZN => n2798);
   U1851 : AOI22_X1 port map( A1 => n2801, A2 => n2800, B1 => n2799, B2 => 
                           n2798, ZN => n2802);
   U1852 : OAI221_X1 port map( B1 => n2806, B2 => n2805, C1 => n2804, C2 => 
                           n2803, A => n2802, ZN => N96);
   U1853 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => n2811, S => n64, Z 
                           => n2166);
   U1854 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => n2813, S => n64, Z 
                           => n2165);
   U1855 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => n2814, S => n64, Z 
                           => n2164);
   U1856 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => n2815, S => n64, Z 
                           => n2163);
   U1857 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => n2816, S => n64, Z 
                           => n2162);
   U1858 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => n2817, S => n64, Z 
                           => n2161);
   U1859 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => n2818, S => n64, Z 
                           => n2160);
   U1860 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => n2819, S => n64, Z 
                           => n2159);
   U1861 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => n2820, S => n64, Z 
                           => n2158);
   U1862 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => n2821, S => n64, Z 
                           => n2157);
   U1863 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => n2822, S => n64, Z 
                           => n2156);
   U1864 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => n2823, S => n64, Z 
                           => n2155);
   U1865 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => n2824, S => n64, Z 
                           => n2154);
   U1866 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => n2825, S => n64, Z 
                           => n2153);
   U1867 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => n2826, S => n64, Z 
                           => n2152);
   U1868 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => n2827, S => n64, Z 
                           => n2151);
   U1869 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => n2828, S => n64, Z 
                           => n2150);
   U1870 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => n2829, S => n64, Z 
                           => n2149);
   U1871 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => n2830, S => n64, Z 
                           => n2148);
   U1872 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => n2831, S => n64, Z 
                           => n2147);
   U1873 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => n2832, S => n64, Z 
                           => n2146);
   U1874 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => n2833, S => n64, Z 
                           => n2145);
   U1875 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => n2834, S => n64, Z 
                           => n2144);
   U1876 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => n2835, S => n64, Z 
                           => n2143);
   U1877 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => n2836, S => n64, Z 
                           => n2142);
   U1878 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => n2837, S => n64, Z 
                           => n2141);
   U1879 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => n2838, S => n64, Z 
                           => n2140);
   U1880 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => n2839, S => n64, Z 
                           => n2139);
   U1881 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => n2840, S => n64, Z 
                           => n2138);
   U1882 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => n2841, S => n64, Z 
                           => n2137);
   U1883 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => n2842, S => n64, Z 
                           => n2136);
   U1884 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => n2843, S => n64, Z 
                           => n2135);
   U1885 : OAI21_X1 port map( B1 => n2844, B2 => n2845, A => n274, ZN => n2812)
                           ;
   U1886 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => n2811, S => 
                           n60_port, Z => n2134);
   U1887 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => n2813, S => 
                           n60_port, Z => n2133);
   U1888 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => n2814, S => 
                           n60_port, Z => n2132);
   U1889 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => n2815, S => 
                           n60_port, Z => n2131);
   U1890 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => n2816, S => 
                           n60_port, Z => n2130);
   U1891 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => n2817, S => 
                           n60_port, Z => n2129);
   U1892 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => n2818, S => 
                           n60_port, Z => n2128);
   U1893 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => n2819, S => 
                           n60_port, Z => n2127);
   U1894 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => n2820, S => 
                           n60_port, Z => n2126);
   U1895 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => n2821, S => 
                           n60_port, Z => n2125);
   U1896 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => n2822, S => 
                           n60_port, Z => n2124);
   U1897 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => n2823, S => 
                           n60_port, Z => n2123);
   U1898 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => n2824, S => 
                           n60_port, Z => n2122);
   U1899 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => n2825, S => 
                           n60_port, Z => n2121);
   U1900 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => n2826, S => 
                           n60_port, Z => n2120);
   U1901 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => n2827, S => 
                           n60_port, Z => n2119);
   U1902 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => n2828, S => 
                           n60_port, Z => n2118);
   U1903 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => n2829, S => 
                           n60_port, Z => n2117);
   U1904 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => n2830, S => 
                           n60_port, Z => n2116);
   U1905 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => n2831, S => 
                           n60_port, Z => n2115);
   U1906 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => n2832, S => 
                           n60_port, Z => n2114);
   U1907 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => n2833, S => 
                           n60_port, Z => n2113);
   U1908 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => n2834, S => n60_port
                           , Z => n2112);
   U1909 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => n2835, S => n60_port
                           , Z => n2111);
   U1910 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => n2836, S => n60_port
                           , Z => n2110);
   U1911 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => n2837, S => n60_port
                           , Z => n2109);
   U1912 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => n2838, S => n60_port
                           , Z => n2108);
   U1913 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => n2839, S => n60_port
                           , Z => n2107);
   U1914 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => n2840, S => n60_port
                           , Z => n2106);
   U1915 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => n2841, S => n60_port
                           , Z => n2105);
   U1916 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => n2842, S => n60_port
                           , Z => n2104);
   U1917 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => n2843, S => n60_port
                           , Z => n2103);
   U1918 : OAI21_X1 port map( B1 => n2844, B2 => n2847, A => n273, ZN => n2846)
                           ;
   U1919 : MUX2_X1 port map( A => REGISTERS_2_31_port, B => n2811, S => 
                           n62_port, Z => n2102);
   U1920 : MUX2_X1 port map( A => REGISTERS_2_30_port, B => n2813, S => 
                           n62_port, Z => n2101);
   U1921 : MUX2_X1 port map( A => REGISTERS_2_29_port, B => n2814, S => 
                           n62_port, Z => n2100);
   U1922 : MUX2_X1 port map( A => REGISTERS_2_28_port, B => n2815, S => 
                           n62_port, Z => n2099);
   U1923 : MUX2_X1 port map( A => REGISTERS_2_27_port, B => n2816, S => 
                           n62_port, Z => n2098);
   U1924 : MUX2_X1 port map( A => REGISTERS_2_26_port, B => n2817, S => 
                           n62_port, Z => n2097);
   U1925 : MUX2_X1 port map( A => REGISTERS_2_25_port, B => n2818, S => 
                           n62_port, Z => n2096);
   U1926 : MUX2_X1 port map( A => REGISTERS_2_24_port, B => n2819, S => 
                           n62_port, Z => n2095);
   U1927 : MUX2_X1 port map( A => REGISTERS_2_23_port, B => n2820, S => 
                           n62_port, Z => n2094);
   U1928 : MUX2_X1 port map( A => REGISTERS_2_22_port, B => n2821, S => 
                           n62_port, Z => n2093);
   U1929 : MUX2_X1 port map( A => REGISTERS_2_21_port, B => n2822, S => 
                           n62_port, Z => n2092);
   U1930 : MUX2_X1 port map( A => REGISTERS_2_20_port, B => n2823, S => 
                           n62_port, Z => n2091);
   U1931 : MUX2_X1 port map( A => REGISTERS_2_19_port, B => n2824, S => 
                           n62_port, Z => n2090);
   U1932 : MUX2_X1 port map( A => REGISTERS_2_18_port, B => n2825, S => 
                           n62_port, Z => n2089);
   U1933 : MUX2_X1 port map( A => REGISTERS_2_17_port, B => n2826, S => 
                           n62_port, Z => n2088);
   U1934 : MUX2_X1 port map( A => REGISTERS_2_16_port, B => n2827, S => 
                           n62_port, Z => n2087);
   U1935 : MUX2_X1 port map( A => REGISTERS_2_15_port, B => n2828, S => 
                           n62_port, Z => n2086);
   U1936 : MUX2_X1 port map( A => REGISTERS_2_14_port, B => n2829, S => 
                           n62_port, Z => n2085);
   U1937 : MUX2_X1 port map( A => REGISTERS_2_13_port, B => n2830, S => 
                           n62_port, Z => n2084);
   U1938 : MUX2_X1 port map( A => REGISTERS_2_12_port, B => n2831, S => 
                           n62_port, Z => n2083);
   U1939 : MUX2_X1 port map( A => REGISTERS_2_11_port, B => n2832, S => 
                           n62_port, Z => n2082);
   U1940 : MUX2_X1 port map( A => REGISTERS_2_10_port, B => n2833, S => 
                           n62_port, Z => n2081);
   U1941 : MUX2_X1 port map( A => REGISTERS_2_9_port, B => n2834, S => n62_port
                           , Z => n2080);
   U1942 : MUX2_X1 port map( A => REGISTERS_2_8_port, B => n2835, S => n62_port
                           , Z => n2079);
   U1943 : MUX2_X1 port map( A => REGISTERS_2_7_port, B => n2836, S => n62_port
                           , Z => n2078);
   U1944 : MUX2_X1 port map( A => REGISTERS_2_6_port, B => n2837, S => n62_port
                           , Z => n2077);
   U1945 : MUX2_X1 port map( A => REGISTERS_2_5_port, B => n2838, S => n62_port
                           , Z => n2076);
   U1946 : MUX2_X1 port map( A => REGISTERS_2_4_port, B => n2839, S => n62_port
                           , Z => n2075);
   U1947 : MUX2_X1 port map( A => REGISTERS_2_3_port, B => n2840, S => n62_port
                           , Z => n2074);
   U1948 : MUX2_X1 port map( A => REGISTERS_2_2_port, B => n2841, S => n62_port
                           , Z => n2073);
   U1949 : MUX2_X1 port map( A => REGISTERS_2_1_port, B => n2842, S => n62_port
                           , Z => n2072);
   U1950 : MUX2_X1 port map( A => REGISTERS_2_0_port, B => n2843, S => n62_port
                           , Z => n2071);
   U1951 : OAI21_X1 port map( B1 => n2844, B2 => n2849, A => n273, ZN => n2848)
                           ;
   U1952 : MUX2_X1 port map( A => REGISTERS_3_31_port, B => n2811, S => 
                           n56_port, Z => n2070);
   U1953 : MUX2_X1 port map( A => REGISTERS_3_30_port, B => n2813, S => 
                           n56_port, Z => n2069);
   U1954 : MUX2_X1 port map( A => REGISTERS_3_29_port, B => n2814, S => 
                           n56_port, Z => n2068);
   U1955 : MUX2_X1 port map( A => REGISTERS_3_28_port, B => n2815, S => 
                           n56_port, Z => n2067);
   U1956 : MUX2_X1 port map( A => REGISTERS_3_27_port, B => n2816, S => 
                           n56_port, Z => n2066);
   U1957 : MUX2_X1 port map( A => REGISTERS_3_26_port, B => n2817, S => 
                           n56_port, Z => n2065);
   U1958 : MUX2_X1 port map( A => REGISTERS_3_25_port, B => n2818, S => 
                           n56_port, Z => n2064);
   U1959 : MUX2_X1 port map( A => REGISTERS_3_24_port, B => n2819, S => 
                           n56_port, Z => n2063);
   U1960 : MUX2_X1 port map( A => REGISTERS_3_23_port, B => n2820, S => 
                           n56_port, Z => n2062);
   U1961 : MUX2_X1 port map( A => REGISTERS_3_22_port, B => n2821, S => 
                           n56_port, Z => n2061);
   U1962 : MUX2_X1 port map( A => REGISTERS_3_21_port, B => n2822, S => 
                           n56_port, Z => n2060);
   U1963 : MUX2_X1 port map( A => REGISTERS_3_20_port, B => n2823, S => 
                           n56_port, Z => n2059);
   U1964 : MUX2_X1 port map( A => REGISTERS_3_19_port, B => n2824, S => 
                           n56_port, Z => n2058);
   U1965 : MUX2_X1 port map( A => REGISTERS_3_18_port, B => n2825, S => 
                           n56_port, Z => n2057);
   U1966 : MUX2_X1 port map( A => REGISTERS_3_17_port, B => n2826, S => 
                           n56_port, Z => n2056);
   U1967 : MUX2_X1 port map( A => REGISTERS_3_16_port, B => n2827, S => 
                           n56_port, Z => n2055);
   U1968 : MUX2_X1 port map( A => REGISTERS_3_15_port, B => n2828, S => 
                           n56_port, Z => n2054);
   U1969 : MUX2_X1 port map( A => REGISTERS_3_14_port, B => n2829, S => 
                           n56_port, Z => n2053);
   U1970 : MUX2_X1 port map( A => REGISTERS_3_13_port, B => n2830, S => 
                           n56_port, Z => n2052);
   U1971 : MUX2_X1 port map( A => REGISTERS_3_12_port, B => n2831, S => 
                           n56_port, Z => n2051);
   U1972 : MUX2_X1 port map( A => REGISTERS_3_11_port, B => n2832, S => 
                           n56_port, Z => n2050);
   U1973 : MUX2_X1 port map( A => REGISTERS_3_10_port, B => n2833, S => 
                           n56_port, Z => n2049);
   U1974 : MUX2_X1 port map( A => REGISTERS_3_9_port, B => n2834, S => n56_port
                           , Z => n2048);
   U1975 : MUX2_X1 port map( A => REGISTERS_3_8_port, B => n2835, S => n56_port
                           , Z => n2047);
   U1976 : MUX2_X1 port map( A => REGISTERS_3_7_port, B => n2836, S => n56_port
                           , Z => n2046);
   U1977 : MUX2_X1 port map( A => REGISTERS_3_6_port, B => n2837, S => n56_port
                           , Z => n2045);
   U1978 : MUX2_X1 port map( A => REGISTERS_3_5_port, B => n2838, S => n56_port
                           , Z => n2044);
   U1979 : MUX2_X1 port map( A => REGISTERS_3_4_port, B => n2839, S => n56_port
                           , Z => n2043);
   U1980 : MUX2_X1 port map( A => REGISTERS_3_3_port, B => n2840, S => n56_port
                           , Z => n2042);
   U1981 : MUX2_X1 port map( A => REGISTERS_3_2_port, B => n2841, S => n56_port
                           , Z => n2041);
   U1982 : MUX2_X1 port map( A => REGISTERS_3_1_port, B => n2842, S => n56_port
                           , Z => n2040);
   U1983 : MUX2_X1 port map( A => REGISTERS_3_0_port, B => n2843, S => n56_port
                           , Z => n2039);
   U1984 : OAI21_X1 port map( B1 => n2844, B2 => n2851, A => n273, ZN => n2850)
                           ;
   U1985 : MUX2_X1 port map( A => REGISTERS_4_31_port, B => n2811, S => 
                           n58_port, Z => n2038);
   U1986 : MUX2_X1 port map( A => REGISTERS_4_30_port, B => n2813, S => 
                           n58_port, Z => n2037);
   U1987 : MUX2_X1 port map( A => REGISTERS_4_29_port, B => n2814, S => 
                           n58_port, Z => n2036);
   U1988 : MUX2_X1 port map( A => REGISTERS_4_28_port, B => n2815, S => 
                           n58_port, Z => n2035);
   U1989 : MUX2_X1 port map( A => REGISTERS_4_27_port, B => n2816, S => 
                           n58_port, Z => n2034);
   U1990 : MUX2_X1 port map( A => REGISTERS_4_26_port, B => n2817, S => 
                           n58_port, Z => n2033);
   U1991 : MUX2_X1 port map( A => REGISTERS_4_25_port, B => n2818, S => 
                           n58_port, Z => n2032);
   U1992 : MUX2_X1 port map( A => REGISTERS_4_24_port, B => n2819, S => 
                           n58_port, Z => n2031);
   U1993 : MUX2_X1 port map( A => REGISTERS_4_23_port, B => n2820, S => 
                           n58_port, Z => n2030);
   U1994 : MUX2_X1 port map( A => REGISTERS_4_22_port, B => n2821, S => 
                           n58_port, Z => n2029);
   U1995 : MUX2_X1 port map( A => REGISTERS_4_21_port, B => n2822, S => 
                           n58_port, Z => n2028);
   U1996 : MUX2_X1 port map( A => REGISTERS_4_20_port, B => n2823, S => 
                           n58_port, Z => n2027);
   U1997 : MUX2_X1 port map( A => REGISTERS_4_19_port, B => n2824, S => 
                           n58_port, Z => n2026);
   U1998 : MUX2_X1 port map( A => REGISTERS_4_18_port, B => n2825, S => 
                           n58_port, Z => n2025);
   U1999 : MUX2_X1 port map( A => REGISTERS_4_17_port, B => n2826, S => 
                           n58_port, Z => n2024);
   U2000 : MUX2_X1 port map( A => REGISTERS_4_16_port, B => n2827, S => 
                           n58_port, Z => n2023);
   U2001 : MUX2_X1 port map( A => REGISTERS_4_15_port, B => n2828, S => 
                           n58_port, Z => n2022);
   U2002 : MUX2_X1 port map( A => REGISTERS_4_14_port, B => n2829, S => 
                           n58_port, Z => n2021);
   U2003 : MUX2_X1 port map( A => REGISTERS_4_13_port, B => n2830, S => 
                           n58_port, Z => n2020);
   U2004 : MUX2_X1 port map( A => REGISTERS_4_12_port, B => n2831, S => 
                           n58_port, Z => n2019);
   U2005 : MUX2_X1 port map( A => REGISTERS_4_11_port, B => n2832, S => 
                           n58_port, Z => n2018);
   U2006 : MUX2_X1 port map( A => REGISTERS_4_10_port, B => n2833, S => 
                           n58_port, Z => n2017);
   U2007 : MUX2_X1 port map( A => REGISTERS_4_9_port, B => n2834, S => n58_port
                           , Z => n2016);
   U2008 : MUX2_X1 port map( A => REGISTERS_4_8_port, B => n2835, S => n58_port
                           , Z => n2015);
   U2009 : MUX2_X1 port map( A => REGISTERS_4_7_port, B => n2836, S => n58_port
                           , Z => n2014);
   U2010 : MUX2_X1 port map( A => REGISTERS_4_6_port, B => n2837, S => n58_port
                           , Z => n2013);
   U2011 : MUX2_X1 port map( A => REGISTERS_4_5_port, B => n2838, S => n58_port
                           , Z => n2012);
   U2012 : MUX2_X1 port map( A => REGISTERS_4_4_port, B => n2839, S => n58_port
                           , Z => n2011);
   U2013 : MUX2_X1 port map( A => REGISTERS_4_3_port, B => n2840, S => n58_port
                           , Z => n2010);
   U2014 : MUX2_X1 port map( A => REGISTERS_4_2_port, B => n2841, S => n58_port
                           , Z => n2009);
   U2015 : MUX2_X1 port map( A => REGISTERS_4_1_port, B => n2842, S => n58_port
                           , Z => n2008);
   U2016 : MUX2_X1 port map( A => REGISTERS_4_0_port, B => n2843, S => n58_port
                           , Z => n2007);
   U2017 : OAI21_X1 port map( B1 => n2844, B2 => n2853, A => n273, ZN => n2852)
                           ;
   U2018 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => n2811, S => 
                           n52_port, Z => n2006);
   U2019 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => n2813, S => 
                           n52_port, Z => n2005);
   U2020 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => n2814, S => 
                           n52_port, Z => n2004);
   U2021 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => n2815, S => 
                           n52_port, Z => n2003);
   U2022 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => n2816, S => 
                           n52_port, Z => n2002);
   U2023 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => n2817, S => 
                           n52_port, Z => n2001);
   U2024 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => n2818, S => 
                           n52_port, Z => n2000);
   U2025 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => n2819, S => 
                           n52_port, Z => n1999);
   U2026 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => n2820, S => 
                           n52_port, Z => n1998);
   U2027 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => n2821, S => 
                           n52_port, Z => n1997);
   U2028 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => n2822, S => 
                           n52_port, Z => n1996);
   U2029 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => n2823, S => 
                           n52_port, Z => n1995);
   U2030 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => n2824, S => 
                           n52_port, Z => n1994);
   U2031 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => n2825, S => 
                           n52_port, Z => n1993);
   U2032 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => n2826, S => 
                           n52_port, Z => n1992);
   U2033 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => n2827, S => 
                           n52_port, Z => n1991);
   U2034 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => n2828, S => 
                           n52_port, Z => n1990);
   U2035 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => n2829, S => 
                           n52_port, Z => n1989);
   U2036 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => n2830, S => 
                           n52_port, Z => n1988);
   U2037 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => n2831, S => 
                           n52_port, Z => n1987);
   U2038 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => n2832, S => 
                           n52_port, Z => n1986);
   U2039 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => n2833, S => 
                           n52_port, Z => n1985);
   U2040 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => n2834, S => n52_port
                           , Z => n1984);
   U2041 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => n2835, S => n52_port
                           , Z => n1983);
   U2042 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => n2836, S => n52_port
                           , Z => n1982);
   U2043 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => n2837, S => n52_port
                           , Z => n1981);
   U2044 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => n2838, S => n52_port
                           , Z => n1980);
   U2045 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => n2839, S => n52_port
                           , Z => n1979);
   U2046 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => n2840, S => n52_port
                           , Z => n1978);
   U2047 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => n2841, S => n52_port
                           , Z => n1977);
   U2048 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => n2842, S => n52_port
                           , Z => n1976);
   U2049 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => n2843, S => n52_port
                           , Z => n1975);
   U2050 : OAI21_X1 port map( B1 => n2844, B2 => n2855, A => n273, ZN => n2854)
                           ;
   U2051 : MUX2_X1 port map( A => REGISTERS_6_31_port, B => n2811, S => 
                           n54_port, Z => n1974);
   U2052 : MUX2_X1 port map( A => REGISTERS_6_30_port, B => n2813, S => 
                           n54_port, Z => n1973);
   U2053 : MUX2_X1 port map( A => REGISTERS_6_29_port, B => n2814, S => 
                           n54_port, Z => n1972);
   U2054 : MUX2_X1 port map( A => REGISTERS_6_28_port, B => n2815, S => 
                           n54_port, Z => n1971);
   U2055 : MUX2_X1 port map( A => REGISTERS_6_27_port, B => n2816, S => 
                           n54_port, Z => n1970);
   U2056 : MUX2_X1 port map( A => REGISTERS_6_26_port, B => n2817, S => 
                           n54_port, Z => n1969);
   U2057 : MUX2_X1 port map( A => REGISTERS_6_25_port, B => n2818, S => 
                           n54_port, Z => n1968);
   U2058 : MUX2_X1 port map( A => REGISTERS_6_24_port, B => n2819, S => 
                           n54_port, Z => n1967);
   U2059 : MUX2_X1 port map( A => REGISTERS_6_23_port, B => n2820, S => 
                           n54_port, Z => n1966);
   U2060 : MUX2_X1 port map( A => REGISTERS_6_22_port, B => n2821, S => 
                           n54_port, Z => n1965);
   U2061 : MUX2_X1 port map( A => REGISTERS_6_21_port, B => n2822, S => 
                           n54_port, Z => n1964);
   U2062 : MUX2_X1 port map( A => REGISTERS_6_20_port, B => n2823, S => 
                           n54_port, Z => n1963);
   U2063 : MUX2_X1 port map( A => REGISTERS_6_19_port, B => n2824, S => 
                           n54_port, Z => n1962);
   U2064 : MUX2_X1 port map( A => REGISTERS_6_18_port, B => n2825, S => 
                           n54_port, Z => n1961);
   U2065 : MUX2_X1 port map( A => REGISTERS_6_17_port, B => n2826, S => 
                           n54_port, Z => n1960);
   U2066 : MUX2_X1 port map( A => REGISTERS_6_16_port, B => n2827, S => 
                           n54_port, Z => n1959);
   U2067 : MUX2_X1 port map( A => REGISTERS_6_15_port, B => n2828, S => 
                           n54_port, Z => n1958);
   U2068 : MUX2_X1 port map( A => REGISTERS_6_14_port, B => n2829, S => 
                           n54_port, Z => n1957);
   U2069 : MUX2_X1 port map( A => REGISTERS_6_13_port, B => n2830, S => 
                           n54_port, Z => n1956);
   U2070 : MUX2_X1 port map( A => REGISTERS_6_12_port, B => n2831, S => 
                           n54_port, Z => n1955);
   U2071 : MUX2_X1 port map( A => REGISTERS_6_11_port, B => n2832, S => 
                           n54_port, Z => n1954);
   U2072 : MUX2_X1 port map( A => REGISTERS_6_10_port, B => n2833, S => 
                           n54_port, Z => n1953);
   U2073 : MUX2_X1 port map( A => REGISTERS_6_9_port, B => n2834, S => n54_port
                           , Z => n1952);
   U2074 : MUX2_X1 port map( A => REGISTERS_6_8_port, B => n2835, S => n54_port
                           , Z => n1951);
   U2075 : MUX2_X1 port map( A => REGISTERS_6_7_port, B => n2836, S => n54_port
                           , Z => n1950);
   U2076 : MUX2_X1 port map( A => REGISTERS_6_6_port, B => n2837, S => n54_port
                           , Z => n1949);
   U2077 : MUX2_X1 port map( A => REGISTERS_6_5_port, B => n2838, S => n54_port
                           , Z => n1948);
   U2078 : MUX2_X1 port map( A => REGISTERS_6_4_port, B => n2839, S => n54_port
                           , Z => n1947);
   U2079 : MUX2_X1 port map( A => REGISTERS_6_3_port, B => n2840, S => n54_port
                           , Z => n1946);
   U2080 : MUX2_X1 port map( A => REGISTERS_6_2_port, B => n2841, S => n54_port
                           , Z => n1945);
   U2081 : MUX2_X1 port map( A => REGISTERS_6_1_port, B => n2842, S => n54_port
                           , Z => n1944);
   U2082 : MUX2_X1 port map( A => REGISTERS_6_0_port, B => n2843, S => n54_port
                           , Z => n1943);
   U2083 : OAI21_X1 port map( B1 => n2844, B2 => n2857, A => n273, ZN => n2856)
                           ;
   U2084 : MUX2_X1 port map( A => REGISTERS_7_31_port, B => n2811, S => 
                           n48_port, Z => n1942);
   U2085 : MUX2_X1 port map( A => REGISTERS_7_30_port, B => n2813, S => 
                           n48_port, Z => n1941);
   U2086 : MUX2_X1 port map( A => REGISTERS_7_29_port, B => n2814, S => 
                           n48_port, Z => n1940);
   U2087 : MUX2_X1 port map( A => REGISTERS_7_28_port, B => n2815, S => 
                           n48_port, Z => n1939);
   U2088 : MUX2_X1 port map( A => REGISTERS_7_27_port, B => n2816, S => 
                           n48_port, Z => n1938);
   U2089 : MUX2_X1 port map( A => REGISTERS_7_26_port, B => n2817, S => 
                           n48_port, Z => n1937);
   U2090 : MUX2_X1 port map( A => REGISTERS_7_25_port, B => n2818, S => 
                           n48_port, Z => n1936);
   U2091 : MUX2_X1 port map( A => REGISTERS_7_24_port, B => n2819, S => 
                           n48_port, Z => n1935);
   U2092 : MUX2_X1 port map( A => REGISTERS_7_23_port, B => n2820, S => 
                           n48_port, Z => n1934);
   U2093 : MUX2_X1 port map( A => REGISTERS_7_22_port, B => n2821, S => 
                           n48_port, Z => n1933);
   U2094 : MUX2_X1 port map( A => REGISTERS_7_21_port, B => n2822, S => 
                           n48_port, Z => n1932);
   U2095 : MUX2_X1 port map( A => REGISTERS_7_20_port, B => n2823, S => 
                           n48_port, Z => n1931);
   U2096 : MUX2_X1 port map( A => REGISTERS_7_19_port, B => n2824, S => 
                           n48_port, Z => n1930);
   U2097 : MUX2_X1 port map( A => REGISTERS_7_18_port, B => n2825, S => 
                           n48_port, Z => n1929);
   U2098 : MUX2_X1 port map( A => REGISTERS_7_17_port, B => n2826, S => 
                           n48_port, Z => n1928);
   U2099 : MUX2_X1 port map( A => REGISTERS_7_16_port, B => n2827, S => 
                           n48_port, Z => n1927);
   U2100 : MUX2_X1 port map( A => REGISTERS_7_15_port, B => n2828, S => 
                           n48_port, Z => n1926);
   U2101 : MUX2_X1 port map( A => REGISTERS_7_14_port, B => n2829, S => 
                           n48_port, Z => n1925);
   U2102 : MUX2_X1 port map( A => REGISTERS_7_13_port, B => n2830, S => 
                           n48_port, Z => n1924);
   U2103 : MUX2_X1 port map( A => REGISTERS_7_12_port, B => n2831, S => 
                           n48_port, Z => n1923);
   U2104 : MUX2_X1 port map( A => REGISTERS_7_11_port, B => n2832, S => 
                           n48_port, Z => n1922);
   U2105 : MUX2_X1 port map( A => REGISTERS_7_10_port, B => n2833, S => 
                           n48_port, Z => n1921);
   U2106 : MUX2_X1 port map( A => REGISTERS_7_9_port, B => n2834, S => n48_port
                           , Z => n1920);
   U2107 : MUX2_X1 port map( A => REGISTERS_7_8_port, B => n2835, S => n48_port
                           , Z => n1919);
   U2108 : MUX2_X1 port map( A => REGISTERS_7_7_port, B => n2836, S => n48_port
                           , Z => n1918);
   U2109 : MUX2_X1 port map( A => REGISTERS_7_6_port, B => n2837, S => n48_port
                           , Z => n1917);
   U2110 : MUX2_X1 port map( A => REGISTERS_7_5_port, B => n2838, S => n48_port
                           , Z => n1916);
   U2111 : MUX2_X1 port map( A => REGISTERS_7_4_port, B => n2839, S => n48_port
                           , Z => n1915);
   U2112 : MUX2_X1 port map( A => REGISTERS_7_3_port, B => n2840, S => n48_port
                           , Z => n1914);
   U2113 : MUX2_X1 port map( A => REGISTERS_7_2_port, B => n2841, S => n48_port
                           , Z => n1913);
   U2114 : MUX2_X1 port map( A => REGISTERS_7_1_port, B => n2842, S => n48_port
                           , Z => n1912);
   U2115 : MUX2_X1 port map( A => REGISTERS_7_0_port, B => n2843, S => n48_port
                           , Z => n1911);
   U2116 : OAI21_X1 port map( B1 => n2844, B2 => n2859, A => n273, ZN => n2858)
                           ;
   U2117 : NAND3_X1 port map( A1 => n2860, A2 => n2861, A3 => n2862, ZN => 
                           n2844);
   U2118 : MUX2_X1 port map( A => REGISTERS_8_31_port, B => n2811, S => 
                           n50_port, Z => n1910);
   U2119 : MUX2_X1 port map( A => REGISTERS_8_30_port, B => n2813, S => 
                           n50_port, Z => n1909);
   U2120 : MUX2_X1 port map( A => REGISTERS_8_29_port, B => n2814, S => 
                           n50_port, Z => n1908);
   U2121 : MUX2_X1 port map( A => REGISTERS_8_28_port, B => n2815, S => 
                           n50_port, Z => n1907);
   U2122 : MUX2_X1 port map( A => REGISTERS_8_27_port, B => n2816, S => 
                           n50_port, Z => n1906);
   U2123 : MUX2_X1 port map( A => REGISTERS_8_26_port, B => n2817, S => 
                           n50_port, Z => n1905);
   U2124 : MUX2_X1 port map( A => REGISTERS_8_25_port, B => n2818, S => 
                           n50_port, Z => n1904);
   U2125 : MUX2_X1 port map( A => REGISTERS_8_24_port, B => n2819, S => 
                           n50_port, Z => n1903);
   U2126 : MUX2_X1 port map( A => REGISTERS_8_23_port, B => n2820, S => 
                           n50_port, Z => n1902);
   U2127 : MUX2_X1 port map( A => REGISTERS_8_22_port, B => n2821, S => 
                           n50_port, Z => n1901);
   U2128 : MUX2_X1 port map( A => REGISTERS_8_21_port, B => n2822, S => 
                           n50_port, Z => n1900);
   U2129 : MUX2_X1 port map( A => REGISTERS_8_20_port, B => n2823, S => 
                           n50_port, Z => n1899);
   U2130 : MUX2_X1 port map( A => REGISTERS_8_19_port, B => n2824, S => 
                           n50_port, Z => n1898);
   U2131 : MUX2_X1 port map( A => REGISTERS_8_18_port, B => n2825, S => 
                           n50_port, Z => n1897);
   U2132 : MUX2_X1 port map( A => REGISTERS_8_17_port, B => n2826, S => 
                           n50_port, Z => n1896);
   U2133 : MUX2_X1 port map( A => REGISTERS_8_16_port, B => n2827, S => 
                           n50_port, Z => n1895);
   U2134 : MUX2_X1 port map( A => REGISTERS_8_15_port, B => n2828, S => 
                           n50_port, Z => n1894);
   U2135 : MUX2_X1 port map( A => REGISTERS_8_14_port, B => n2829, S => 
                           n50_port, Z => n1893);
   U2136 : MUX2_X1 port map( A => REGISTERS_8_13_port, B => n2830, S => 
                           n50_port, Z => n1892);
   U2137 : MUX2_X1 port map( A => REGISTERS_8_12_port, B => n2831, S => 
                           n50_port, Z => n1891);
   U2138 : MUX2_X1 port map( A => REGISTERS_8_11_port, B => n2832, S => 
                           n50_port, Z => n1890);
   U2139 : MUX2_X1 port map( A => REGISTERS_8_10_port, B => n2833, S => 
                           n50_port, Z => n1889);
   U2140 : MUX2_X1 port map( A => REGISTERS_8_9_port, B => n2834, S => n50_port
                           , Z => n1888);
   U2141 : MUX2_X1 port map( A => REGISTERS_8_8_port, B => n2835, S => n50_port
                           , Z => n1887);
   U2142 : MUX2_X1 port map( A => REGISTERS_8_7_port, B => n2836, S => n50_port
                           , Z => n1886);
   U2143 : MUX2_X1 port map( A => REGISTERS_8_6_port, B => n2837, S => n50_port
                           , Z => n1885);
   U2144 : MUX2_X1 port map( A => REGISTERS_8_5_port, B => n2838, S => n50_port
                           , Z => n1884);
   U2145 : MUX2_X1 port map( A => REGISTERS_8_4_port, B => n2839, S => n50_port
                           , Z => n1883);
   U2146 : MUX2_X1 port map( A => REGISTERS_8_3_port, B => n2840, S => n50_port
                           , Z => n1882);
   U2147 : MUX2_X1 port map( A => REGISTERS_8_2_port, B => n2841, S => n50_port
                           , Z => n1881);
   U2148 : MUX2_X1 port map( A => REGISTERS_8_1_port, B => n2842, S => n50_port
                           , Z => n1880);
   U2149 : MUX2_X1 port map( A => REGISTERS_8_0_port, B => n2843, S => n50_port
                           , Z => n1879);
   U2150 : OAI21_X1 port map( B1 => n2845, B2 => n2864, A => n273, ZN => n2863)
                           ;
   U2151 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => n2811, S => 
                           n44_port, Z => n1878);
   U2152 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => n2813, S => 
                           n44_port, Z => n1877);
   U2153 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => n2814, S => 
                           n44_port, Z => n1876);
   U2154 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => n2815, S => 
                           n44_port, Z => n1875);
   U2155 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => n2816, S => 
                           n44_port, Z => n1874);
   U2156 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => n2817, S => 
                           n44_port, Z => n1873);
   U2157 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => n2818, S => 
                           n44_port, Z => n1872);
   U2158 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => n2819, S => 
                           n44_port, Z => n1871);
   U2159 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => n2820, S => 
                           n44_port, Z => n1870);
   U2160 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => n2821, S => 
                           n44_port, Z => n1869);
   U2161 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => n2822, S => 
                           n44_port, Z => n1868);
   U2162 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => n2823, S => 
                           n44_port, Z => n1867);
   U2163 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => n2824, S => 
                           n44_port, Z => n1866);
   U2164 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => n2825, S => 
                           n44_port, Z => n1865);
   U2165 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => n2826, S => 
                           n44_port, Z => n1864);
   U2166 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => n2827, S => 
                           n44_port, Z => n1863);
   U2167 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => n2828, S => 
                           n44_port, Z => n1862);
   U2168 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => n2829, S => 
                           n44_port, Z => n1861);
   U2169 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => n2830, S => 
                           n44_port, Z => n1860);
   U2170 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => n2831, S => 
                           n44_port, Z => n1859);
   U2171 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => n2832, S => 
                           n44_port, Z => n1858);
   U2172 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => n2833, S => 
                           n44_port, Z => n1857);
   U2173 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => n2834, S => n44_port
                           , Z => n1856);
   U2174 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => n2835, S => n44_port
                           , Z => n1855);
   U2175 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => n2836, S => n44_port
                           , Z => n1854);
   U2176 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => n2837, S => n44_port
                           , Z => n1853);
   U2177 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => n2838, S => n44_port
                           , Z => n1852);
   U2178 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => n2839, S => n44_port
                           , Z => n1851);
   U2179 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => n2840, S => n44_port
                           , Z => n1850);
   U2180 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => n2841, S => n44_port
                           , Z => n1849);
   U2181 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => n2842, S => n44_port
                           , Z => n1848);
   U2182 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => n2843, S => n44_port
                           , Z => n1847);
   U2183 : OAI21_X1 port map( B1 => n2847, B2 => n2864, A => n273, ZN => n2865)
                           ;
   U2184 : MUX2_X1 port map( A => REGISTERS_10_31_port, B => n2811, S => 
                           n46_port, Z => n1846);
   U2185 : MUX2_X1 port map( A => REGISTERS_10_30_port, B => n2813, S => 
                           n46_port, Z => n1845);
   U2186 : MUX2_X1 port map( A => REGISTERS_10_29_port, B => n2814, S => 
                           n46_port, Z => n1844);
   U2187 : MUX2_X1 port map( A => REGISTERS_10_28_port, B => n2815, S => 
                           n46_port, Z => n1843);
   U2188 : MUX2_X1 port map( A => REGISTERS_10_27_port, B => n2816, S => 
                           n46_port, Z => n1842);
   U2189 : MUX2_X1 port map( A => REGISTERS_10_26_port, B => n2817, S => 
                           n46_port, Z => n1841);
   U2190 : MUX2_X1 port map( A => REGISTERS_10_25_port, B => n2818, S => 
                           n46_port, Z => n1840);
   U2191 : MUX2_X1 port map( A => REGISTERS_10_24_port, B => n2819, S => 
                           n46_port, Z => n1839);
   U2192 : MUX2_X1 port map( A => REGISTERS_10_23_port, B => n2820, S => 
                           n46_port, Z => n1838);
   U2193 : MUX2_X1 port map( A => REGISTERS_10_22_port, B => n2821, S => 
                           n46_port, Z => n1837);
   U2194 : MUX2_X1 port map( A => REGISTERS_10_21_port, B => n2822, S => 
                           n46_port, Z => n1836);
   U2195 : MUX2_X1 port map( A => REGISTERS_10_20_port, B => n2823, S => 
                           n46_port, Z => n1835);
   U2196 : MUX2_X1 port map( A => REGISTERS_10_19_port, B => n2824, S => 
                           n46_port, Z => n1834);
   U2197 : MUX2_X1 port map( A => REGISTERS_10_18_port, B => n2825, S => 
                           n46_port, Z => n1833);
   U2198 : MUX2_X1 port map( A => REGISTERS_10_17_port, B => n2826, S => 
                           n46_port, Z => n1832);
   U2199 : MUX2_X1 port map( A => REGISTERS_10_16_port, B => n2827, S => 
                           n46_port, Z => n1831);
   U2200 : MUX2_X1 port map( A => REGISTERS_10_15_port, B => n2828, S => 
                           n46_port, Z => n1830);
   U2201 : MUX2_X1 port map( A => REGISTERS_10_14_port, B => n2829, S => 
                           n46_port, Z => n1829);
   U2202 : MUX2_X1 port map( A => REGISTERS_10_13_port, B => n2830, S => 
                           n46_port, Z => n1828);
   U2203 : MUX2_X1 port map( A => REGISTERS_10_12_port, B => n2831, S => 
                           n46_port, Z => n1827);
   U2204 : MUX2_X1 port map( A => REGISTERS_10_11_port, B => n2832, S => 
                           n46_port, Z => n1826);
   U2205 : MUX2_X1 port map( A => REGISTERS_10_10_port, B => n2833, S => 
                           n46_port, Z => n1825);
   U2206 : MUX2_X1 port map( A => REGISTERS_10_9_port, B => n2834, S => 
                           n46_port, Z => n1824);
   U2207 : MUX2_X1 port map( A => REGISTERS_10_8_port, B => n2835, S => 
                           n46_port, Z => n1823);
   U2208 : MUX2_X1 port map( A => REGISTERS_10_7_port, B => n2836, S => 
                           n46_port, Z => n1822);
   U2209 : MUX2_X1 port map( A => REGISTERS_10_6_port, B => n2837, S => 
                           n46_port, Z => n1821);
   U2210 : MUX2_X1 port map( A => REGISTERS_10_5_port, B => n2838, S => 
                           n46_port, Z => n1820);
   U2211 : MUX2_X1 port map( A => REGISTERS_10_4_port, B => n2839, S => 
                           n46_port, Z => n1819);
   U2212 : MUX2_X1 port map( A => REGISTERS_10_3_port, B => n2840, S => 
                           n46_port, Z => n1818);
   U2213 : MUX2_X1 port map( A => REGISTERS_10_2_port, B => n2841, S => 
                           n46_port, Z => n1817);
   U2214 : MUX2_X1 port map( A => REGISTERS_10_1_port, B => n2842, S => 
                           n46_port, Z => n1816);
   U2215 : MUX2_X1 port map( A => REGISTERS_10_0_port, B => n2843, S => 
                           n46_port, Z => n1815);
   U2216 : OAI21_X1 port map( B1 => n2849, B2 => n2864, A => n273, ZN => n2866)
                           ;
   U2217 : MUX2_X1 port map( A => REGISTERS_11_31_port, B => n2811, S => 
                           n40_port, Z => n1814);
   U2218 : MUX2_X1 port map( A => REGISTERS_11_30_port, B => n2813, S => 
                           n40_port, Z => n1813);
   U2219 : MUX2_X1 port map( A => REGISTERS_11_29_port, B => n2814, S => 
                           n40_port, Z => n1812);
   U2220 : MUX2_X1 port map( A => REGISTERS_11_28_port, B => n2815, S => 
                           n40_port, Z => n1811);
   U2221 : MUX2_X1 port map( A => REGISTERS_11_27_port, B => n2816, S => 
                           n40_port, Z => n1810);
   U2222 : MUX2_X1 port map( A => REGISTERS_11_26_port, B => n2817, S => 
                           n40_port, Z => n1809);
   U2223 : MUX2_X1 port map( A => REGISTERS_11_25_port, B => n2818, S => 
                           n40_port, Z => n1808);
   U2224 : MUX2_X1 port map( A => REGISTERS_11_24_port, B => n2819, S => 
                           n40_port, Z => n1807);
   U2225 : MUX2_X1 port map( A => REGISTERS_11_23_port, B => n2820, S => 
                           n40_port, Z => n1806);
   U2226 : MUX2_X1 port map( A => REGISTERS_11_22_port, B => n2821, S => 
                           n40_port, Z => n1805);
   U2227 : MUX2_X1 port map( A => REGISTERS_11_21_port, B => n2822, S => 
                           n40_port, Z => n1804);
   U2228 : MUX2_X1 port map( A => REGISTERS_11_20_port, B => n2823, S => 
                           n40_port, Z => n1803);
   U2229 : MUX2_X1 port map( A => REGISTERS_11_19_port, B => n2824, S => 
                           n40_port, Z => n1802);
   U2230 : MUX2_X1 port map( A => REGISTERS_11_18_port, B => n2825, S => 
                           n40_port, Z => n1801);
   U2231 : MUX2_X1 port map( A => REGISTERS_11_17_port, B => n2826, S => 
                           n40_port, Z => n1800);
   U2232 : MUX2_X1 port map( A => REGISTERS_11_16_port, B => n2827, S => 
                           n40_port, Z => n1799);
   U2233 : MUX2_X1 port map( A => REGISTERS_11_15_port, B => n2828, S => 
                           n40_port, Z => n1798);
   U2234 : MUX2_X1 port map( A => REGISTERS_11_14_port, B => n2829, S => 
                           n40_port, Z => n1797);
   U2235 : MUX2_X1 port map( A => REGISTERS_11_13_port, B => n2830, S => 
                           n40_port, Z => n1796);
   U2236 : MUX2_X1 port map( A => REGISTERS_11_12_port, B => n2831, S => 
                           n40_port, Z => n1795);
   U2237 : MUX2_X1 port map( A => REGISTERS_11_11_port, B => n2832, S => 
                           n40_port, Z => n1794);
   U2238 : MUX2_X1 port map( A => REGISTERS_11_10_port, B => n2833, S => 
                           n40_port, Z => n1793);
   U2239 : MUX2_X1 port map( A => REGISTERS_11_9_port, B => n2834, S => 
                           n40_port, Z => n1792);
   U2240 : MUX2_X1 port map( A => REGISTERS_11_8_port, B => n2835, S => 
                           n40_port, Z => n1791);
   U2241 : MUX2_X1 port map( A => REGISTERS_11_7_port, B => n2836, S => 
                           n40_port, Z => n1790);
   U2242 : MUX2_X1 port map( A => REGISTERS_11_6_port, B => n2837, S => 
                           n40_port, Z => n1789);
   U2243 : MUX2_X1 port map( A => REGISTERS_11_5_port, B => n2838, S => 
                           n40_port, Z => n1788);
   U2244 : MUX2_X1 port map( A => REGISTERS_11_4_port, B => n2839, S => 
                           n40_port, Z => n1787);
   U2245 : MUX2_X1 port map( A => REGISTERS_11_3_port, B => n2840, S => 
                           n40_port, Z => n1786);
   U2246 : MUX2_X1 port map( A => REGISTERS_11_2_port, B => n2841, S => 
                           n40_port, Z => n1785);
   U2247 : MUX2_X1 port map( A => REGISTERS_11_1_port, B => n2842, S => 
                           n40_port, Z => n1784);
   U2248 : MUX2_X1 port map( A => REGISTERS_11_0_port, B => n2843, S => 
                           n40_port, Z => n1783);
   U2249 : OAI21_X1 port map( B1 => n2851, B2 => n2864, A => n273, ZN => n2867)
                           ;
   U2250 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => n2811, S => 
                           n42_port, Z => n1782);
   U2251 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => n2813, S => 
                           n42_port, Z => n1781);
   U2252 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => n2814, S => 
                           n42_port, Z => n1780);
   U2253 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => n2815, S => 
                           n42_port, Z => n1779);
   U2254 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => n2816, S => 
                           n42_port, Z => n1778);
   U2255 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => n2817, S => 
                           n42_port, Z => n1777);
   U2256 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => n2818, S => 
                           n42_port, Z => n1776);
   U2257 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => n2819, S => 
                           n42_port, Z => n1775);
   U2258 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => n2820, S => 
                           n42_port, Z => n1774);
   U2259 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => n2821, S => 
                           n42_port, Z => n1773);
   U2260 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => n2822, S => 
                           n42_port, Z => n1772);
   U2261 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => n2823, S => 
                           n42_port, Z => n1771);
   U2262 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => n2824, S => 
                           n42_port, Z => n1770);
   U2263 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => n2825, S => 
                           n42_port, Z => n1769);
   U2264 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => n2826, S => 
                           n42_port, Z => n1768);
   U2265 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => n2827, S => 
                           n42_port, Z => n1767);
   U2266 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => n2828, S => 
                           n42_port, Z => n1766);
   U2267 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => n2829, S => 
                           n42_port, Z => n1765);
   U2268 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => n2830, S => 
                           n42_port, Z => n1764);
   U2269 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => n2831, S => 
                           n42_port, Z => n1763);
   U2270 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => n2832, S => 
                           n42_port, Z => n1762);
   U2271 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => n2833, S => 
                           n42_port, Z => n1761);
   U2272 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => n2834, S => 
                           n42_port, Z => n1760);
   U2273 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => n2835, S => 
                           n42_port, Z => n1759);
   U2274 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => n2836, S => 
                           n42_port, Z => n1758);
   U2275 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => n2837, S => 
                           n42_port, Z => n1757);
   U2276 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => n2838, S => 
                           n42_port, Z => n1756);
   U2277 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => n2839, S => 
                           n42_port, Z => n1755);
   U2278 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => n2840, S => 
                           n42_port, Z => n1754);
   U2279 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => n2841, S => 
                           n42_port, Z => n1753);
   U2280 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => n2842, S => 
                           n42_port, Z => n1752);
   U2281 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => n2843, S => 
                           n42_port, Z => n1751);
   U2282 : OAI21_X1 port map( B1 => n2853, B2 => n2864, A => n274, ZN => n2868)
                           ;
   U2283 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => n2811, S => n2, Z 
                           => n1750);
   U2284 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => n2813, S => n2, Z 
                           => n1749);
   U2285 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => n2814, S => n2, Z 
                           => n1748);
   U2286 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => n2815, S => n2, Z 
                           => n1747);
   U2287 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => n2816, S => n2, Z 
                           => n1746);
   U2288 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => n2817, S => n2, Z 
                           => n1745);
   U2289 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => n2818, S => n2, Z 
                           => n1744);
   U2290 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => n2819, S => n2, Z 
                           => n1743);
   U2291 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => n2820, S => n2, Z 
                           => n1742);
   U2292 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => n2821, S => n2, Z 
                           => n1741);
   U2293 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => n2822, S => n2, Z 
                           => n1740);
   U2294 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => n2823, S => n2, Z 
                           => n1739);
   U2295 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => n2824, S => n2, Z 
                           => n1738);
   U2296 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => n2825, S => n2, Z 
                           => n1737);
   U2297 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => n2826, S => n2, Z 
                           => n1736);
   U2298 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => n2827, S => n2, Z 
                           => n1735);
   U2299 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => n2828, S => n2, Z 
                           => n1734);
   U2300 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => n2829, S => n2, Z 
                           => n1733);
   U2301 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => n2830, S => n2, Z 
                           => n1732);
   U2302 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => n2831, S => n2, Z 
                           => n1731);
   U2303 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => n2832, S => n2, Z 
                           => n1730);
   U2304 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => n2833, S => n2, Z 
                           => n1729);
   U2305 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => n2834, S => n2, Z 
                           => n1728);
   U2306 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => n2835, S => n2, Z 
                           => n1727);
   U2307 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => n2836, S => n2, Z 
                           => n1726);
   U2308 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => n2837, S => n2, Z 
                           => n1725);
   U2309 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => n2838, S => n2, Z 
                           => n1724);
   U2310 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => n2839, S => n2, Z 
                           => n1723);
   U2311 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => n2840, S => n2, Z 
                           => n1722);
   U2312 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => n2841, S => n2, Z 
                           => n1721);
   U2313 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => n2842, S => n2, Z 
                           => n1720);
   U2314 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => n2843, S => n2, Z 
                           => n1719);
   U2315 : OAI21_X1 port map( B1 => n2855, B2 => n2864, A => n274, ZN => n2869)
                           ;
   U2316 : MUX2_X1 port map( A => REGISTERS_14_31_port, B => n2811, S => n4, Z 
                           => n1718);
   U2317 : MUX2_X1 port map( A => REGISTERS_14_30_port, B => n2813, S => n4, Z 
                           => n1717);
   U2318 : MUX2_X1 port map( A => REGISTERS_14_29_port, B => n2814, S => n4, Z 
                           => n1716);
   U2319 : MUX2_X1 port map( A => REGISTERS_14_28_port, B => n2815, S => n4, Z 
                           => n1715);
   U2320 : MUX2_X1 port map( A => REGISTERS_14_27_port, B => n2816, S => n4, Z 
                           => n1714);
   U2321 : MUX2_X1 port map( A => REGISTERS_14_26_port, B => n2817, S => n4, Z 
                           => n1713);
   U2322 : MUX2_X1 port map( A => REGISTERS_14_25_port, B => n2818, S => n4, Z 
                           => n1712);
   U2323 : MUX2_X1 port map( A => REGISTERS_14_24_port, B => n2819, S => n4, Z 
                           => n1711);
   U2324 : MUX2_X1 port map( A => REGISTERS_14_23_port, B => n2820, S => n4, Z 
                           => n1710);
   U2325 : MUX2_X1 port map( A => REGISTERS_14_22_port, B => n2821, S => n4, Z 
                           => n1709);
   U2326 : MUX2_X1 port map( A => REGISTERS_14_21_port, B => n2822, S => n4, Z 
                           => n1708);
   U2327 : MUX2_X1 port map( A => REGISTERS_14_20_port, B => n2823, S => n4, Z 
                           => n1707);
   U2328 : MUX2_X1 port map( A => REGISTERS_14_19_port, B => n2824, S => n4, Z 
                           => n1706);
   U2329 : MUX2_X1 port map( A => REGISTERS_14_18_port, B => n2825, S => n4, Z 
                           => n1705);
   U2330 : MUX2_X1 port map( A => REGISTERS_14_17_port, B => n2826, S => n4, Z 
                           => n1704);
   U2331 : MUX2_X1 port map( A => REGISTERS_14_16_port, B => n2827, S => n4, Z 
                           => n1703);
   U2332 : MUX2_X1 port map( A => REGISTERS_14_15_port, B => n2828, S => n4, Z 
                           => n1702);
   U2333 : MUX2_X1 port map( A => REGISTERS_14_14_port, B => n2829, S => n4, Z 
                           => n1701);
   U2334 : MUX2_X1 port map( A => REGISTERS_14_13_port, B => n2830, S => n4, Z 
                           => n1700);
   U2335 : MUX2_X1 port map( A => REGISTERS_14_12_port, B => n2831, S => n4, Z 
                           => n1699);
   U2336 : MUX2_X1 port map( A => REGISTERS_14_11_port, B => n2832, S => n4, Z 
                           => n1698);
   U2337 : MUX2_X1 port map( A => REGISTERS_14_10_port, B => n2833, S => n4, Z 
                           => n1697);
   U2338 : MUX2_X1 port map( A => REGISTERS_14_9_port, B => n2834, S => n4, Z 
                           => n1696);
   U2339 : MUX2_X1 port map( A => REGISTERS_14_8_port, B => n2835, S => n4, Z 
                           => n1695);
   U2340 : MUX2_X1 port map( A => REGISTERS_14_7_port, B => n2836, S => n4, Z 
                           => n1694);
   U2341 : MUX2_X1 port map( A => REGISTERS_14_6_port, B => n2837, S => n4, Z 
                           => n1693);
   U2342 : MUX2_X1 port map( A => REGISTERS_14_5_port, B => n2838, S => n4, Z 
                           => n1692);
   U2343 : MUX2_X1 port map( A => REGISTERS_14_4_port, B => n2839, S => n4, Z 
                           => n1691);
   U2344 : MUX2_X1 port map( A => REGISTERS_14_3_port, B => n2840, S => n4, Z 
                           => n1690);
   U2345 : MUX2_X1 port map( A => REGISTERS_14_2_port, B => n2841, S => n4, Z 
                           => n1689);
   U2346 : MUX2_X1 port map( A => REGISTERS_14_1_port, B => n2842, S => n4, Z 
                           => n1688);
   U2347 : MUX2_X1 port map( A => REGISTERS_14_0_port, B => n2843, S => n4, Z 
                           => n1687);
   U2348 : OAI21_X1 port map( B1 => n2857, B2 => n2864, A => n274, ZN => n2870)
                           ;
   U2349 : MUX2_X1 port map( A => REGISTERS_15_31_port, B => n2811, S => n6, Z 
                           => n1686);
   U2350 : MUX2_X1 port map( A => REGISTERS_15_30_port, B => n2813, S => n6, Z 
                           => n1685);
   U2351 : MUX2_X1 port map( A => REGISTERS_15_29_port, B => n2814, S => n6, Z 
                           => n1684);
   U2352 : MUX2_X1 port map( A => REGISTERS_15_28_port, B => n2815, S => n6, Z 
                           => n1683);
   U2353 : MUX2_X1 port map( A => REGISTERS_15_27_port, B => n2816, S => n6, Z 
                           => n1682);
   U2354 : MUX2_X1 port map( A => REGISTERS_15_26_port, B => n2817, S => n6, Z 
                           => n1681);
   U2355 : MUX2_X1 port map( A => REGISTERS_15_25_port, B => n2818, S => n6, Z 
                           => n1680);
   U2356 : MUX2_X1 port map( A => REGISTERS_15_24_port, B => n2819, S => n6, Z 
                           => n1679);
   U2357 : MUX2_X1 port map( A => REGISTERS_15_23_port, B => n2820, S => n6, Z 
                           => n1678);
   U2358 : MUX2_X1 port map( A => REGISTERS_15_22_port, B => n2821, S => n6, Z 
                           => n1677);
   U2359 : MUX2_X1 port map( A => REGISTERS_15_21_port, B => n2822, S => n6, Z 
                           => n1676);
   U2360 : MUX2_X1 port map( A => REGISTERS_15_20_port, B => n2823, S => n6, Z 
                           => n1675);
   U2361 : MUX2_X1 port map( A => REGISTERS_15_19_port, B => n2824, S => n6, Z 
                           => n1674);
   U2362 : MUX2_X1 port map( A => REGISTERS_15_18_port, B => n2825, S => n6, Z 
                           => n1673);
   U2363 : MUX2_X1 port map( A => REGISTERS_15_17_port, B => n2826, S => n6, Z 
                           => n1672);
   U2364 : MUX2_X1 port map( A => REGISTERS_15_16_port, B => n2827, S => n6, Z 
                           => n1671);
   U2365 : MUX2_X1 port map( A => REGISTERS_15_15_port, B => n2828, S => n6, Z 
                           => n1670);
   U2366 : MUX2_X1 port map( A => REGISTERS_15_14_port, B => n2829, S => n6, Z 
                           => n1669);
   U2367 : MUX2_X1 port map( A => REGISTERS_15_13_port, B => n2830, S => n6, Z 
                           => n1668);
   U2368 : MUX2_X1 port map( A => REGISTERS_15_12_port, B => n2831, S => n6, Z 
                           => n1667);
   U2369 : MUX2_X1 port map( A => REGISTERS_15_11_port, B => n2832, S => n6, Z 
                           => n1666);
   U2370 : MUX2_X1 port map( A => REGISTERS_15_10_port, B => n2833, S => n6, Z 
                           => n1665);
   U2371 : MUX2_X1 port map( A => REGISTERS_15_9_port, B => n2834, S => n6, Z 
                           => n1664);
   U2372 : MUX2_X1 port map( A => REGISTERS_15_8_port, B => n2835, S => n6, Z 
                           => n1663);
   U2373 : MUX2_X1 port map( A => REGISTERS_15_7_port, B => n2836, S => n6, Z 
                           => n1662);
   U2374 : MUX2_X1 port map( A => REGISTERS_15_6_port, B => n2837, S => n6, Z 
                           => n1661);
   U2375 : MUX2_X1 port map( A => REGISTERS_15_5_port, B => n2838, S => n6, Z 
                           => n1660);
   U2376 : MUX2_X1 port map( A => REGISTERS_15_4_port, B => n2839, S => n6, Z 
                           => n1659);
   U2377 : MUX2_X1 port map( A => REGISTERS_15_3_port, B => n2840, S => n6, Z 
                           => n1658);
   U2378 : MUX2_X1 port map( A => REGISTERS_15_2_port, B => n2841, S => n6, Z 
                           => n1657);
   U2379 : MUX2_X1 port map( A => REGISTERS_15_1_port, B => n2842, S => n6, Z 
                           => n1656);
   U2380 : MUX2_X1 port map( A => REGISTERS_15_0_port, B => n2843, S => n6, Z 
                           => n1655);
   U2381 : OAI21_X1 port map( B1 => n2859, B2 => n2864, A => n274, ZN => n2871)
                           ;
   U2382 : NAND3_X1 port map( A1 => n2862, A2 => n2861, A3 => ADD_WR(3), ZN => 
                           n2864);
   U2383 : INV_X1 port map( A => ADD_WR(4), ZN => n2861);
   U2384 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => n2811, S => n8, Z 
                           => n1654);
   U2385 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => n2813, S => n8, Z 
                           => n1653);
   U2386 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => n2814, S => n8, Z 
                           => n1652);
   U2387 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => n2815, S => n8, Z 
                           => n1651);
   U2388 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => n2816, S => n8, Z 
                           => n1650);
   U2389 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => n2817, S => n8, Z 
                           => n1649);
   U2390 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => n2818, S => n8, Z 
                           => n1648);
   U2391 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => n2819, S => n8, Z 
                           => n1647);
   U2392 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => n2820, S => n8, Z 
                           => n1646);
   U2393 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => n2821, S => n8, Z 
                           => n1645);
   U2394 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => n2822, S => n8, Z 
                           => n1644);
   U2395 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => n2823, S => n8, Z 
                           => n1643);
   U2396 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => n2824, S => n8, Z 
                           => n1642);
   U2397 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => n2825, S => n8, Z 
                           => n1641);
   U2398 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => n2826, S => n8, Z 
                           => n1640);
   U2399 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => n2827, S => n8, Z 
                           => n1639);
   U2400 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => n2828, S => n8, Z 
                           => n1638);
   U2401 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => n2829, S => n8, Z 
                           => n1637);
   U2402 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => n2830, S => n8, Z 
                           => n1636);
   U2403 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => n2831, S => n8, Z 
                           => n1635);
   U2404 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => n2832, S => n8, Z 
                           => n1634);
   U2405 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => n2833, S => n8, Z 
                           => n1633);
   U2406 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => n2834, S => n8, Z 
                           => n1632);
   U2407 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => n2835, S => n8, Z 
                           => n1631);
   U2408 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => n2836, S => n8, Z 
                           => n1630);
   U2409 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => n2837, S => n8, Z 
                           => n1629);
   U2410 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => n2838, S => n8, Z 
                           => n1628);
   U2411 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => n2839, S => n8, Z 
                           => n1627);
   U2412 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => n2840, S => n8, Z 
                           => n1626);
   U2413 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => n2841, S => n8, Z 
                           => n1625);
   U2414 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => n2842, S => n8, Z 
                           => n1624);
   U2415 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => n2843, S => n8, Z 
                           => n1623);
   U2416 : OAI21_X1 port map( B1 => n2845, B2 => n2873, A => n274, ZN => n2872)
                           ;
   U2417 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => n2811, S => n10, Z
                           => n1622);
   U2418 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => n2813, S => n10, Z
                           => n1621);
   U2419 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => n2814, S => n10, Z
                           => n1620);
   U2420 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => n2815, S => n10, Z
                           => n1619);
   U2421 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => n2816, S => n10, Z
                           => n1618);
   U2422 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => n2817, S => n10, Z
                           => n1617);
   U2423 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => n2818, S => n10, Z
                           => n1616);
   U2424 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => n2819, S => n10, Z
                           => n1615);
   U2425 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => n2820, S => n10, Z
                           => n1614);
   U2426 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => n2821, S => n10, Z
                           => n1613);
   U2427 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => n2822, S => n10, Z
                           => n1612);
   U2428 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => n2823, S => n10, Z
                           => n1611);
   U2429 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => n2824, S => n10, Z
                           => n1610);
   U2430 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => n2825, S => n10, Z
                           => n1609);
   U2431 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => n2826, S => n10, Z
                           => n1608);
   U2432 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => n2827, S => n10, Z
                           => n1607);
   U2433 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => n2828, S => n10, Z
                           => n1606);
   U2434 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => n2829, S => n10, Z
                           => n1605);
   U2435 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => n2830, S => n10, Z
                           => n1604);
   U2436 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => n2831, S => n10, Z
                           => n1603);
   U2437 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => n2832, S => n10, Z
                           => n1602);
   U2438 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => n2833, S => n10, Z
                           => n1601);
   U2439 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => n2834, S => n10, Z 
                           => n1600);
   U2440 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => n2835, S => n10, Z 
                           => n1599);
   U2441 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => n2836, S => n10, Z 
                           => n1598);
   U2442 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => n2837, S => n10, Z 
                           => n1597);
   U2443 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => n2838, S => n10, Z 
                           => n1596);
   U2444 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => n2839, S => n10, Z 
                           => n1595);
   U2445 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => n2840, S => n10, Z 
                           => n1594);
   U2446 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => n2841, S => n10, Z 
                           => n1593);
   U2447 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => n2842, S => n10, Z 
                           => n1592);
   U2448 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => n2843, S => n10, Z 
                           => n1591);
   U2449 : OAI21_X1 port map( B1 => n2847, B2 => n2873, A => n274, ZN => n2874)
                           ;
   U2450 : MUX2_X1 port map( A => REGISTERS_18_31_port, B => n2811, S => n12, Z
                           => n1590);
   U2451 : MUX2_X1 port map( A => REGISTERS_18_30_port, B => n2813, S => n12, Z
                           => n1589);
   U2452 : MUX2_X1 port map( A => REGISTERS_18_29_port, B => n2814, S => n12, Z
                           => n1588);
   U2453 : MUX2_X1 port map( A => REGISTERS_18_28_port, B => n2815, S => n12, Z
                           => n1587);
   U2454 : MUX2_X1 port map( A => REGISTERS_18_27_port, B => n2816, S => n12, Z
                           => n1586);
   U2455 : MUX2_X1 port map( A => REGISTERS_18_26_port, B => n2817, S => n12, Z
                           => n1585);
   U2456 : MUX2_X1 port map( A => REGISTERS_18_25_port, B => n2818, S => n12, Z
                           => n1584);
   U2457 : MUX2_X1 port map( A => REGISTERS_18_24_port, B => n2819, S => n12, Z
                           => n1583);
   U2458 : MUX2_X1 port map( A => REGISTERS_18_23_port, B => n2820, S => n12, Z
                           => n1582);
   U2459 : MUX2_X1 port map( A => REGISTERS_18_22_port, B => n2821, S => n12, Z
                           => n1581);
   U2460 : MUX2_X1 port map( A => REGISTERS_18_21_port, B => n2822, S => n12, Z
                           => n1580);
   U2461 : MUX2_X1 port map( A => REGISTERS_18_20_port, B => n2823, S => n12, Z
                           => n1579);
   U2462 : MUX2_X1 port map( A => REGISTERS_18_19_port, B => n2824, S => n12, Z
                           => n1578);
   U2463 : MUX2_X1 port map( A => REGISTERS_18_18_port, B => n2825, S => n12, Z
                           => n1577);
   U2464 : MUX2_X1 port map( A => REGISTERS_18_17_port, B => n2826, S => n12, Z
                           => n1576);
   U2465 : MUX2_X1 port map( A => REGISTERS_18_16_port, B => n2827, S => n12, Z
                           => n1575);
   U2466 : MUX2_X1 port map( A => REGISTERS_18_15_port, B => n2828, S => n12, Z
                           => n1574);
   U2467 : MUX2_X1 port map( A => REGISTERS_18_14_port, B => n2829, S => n12, Z
                           => n1573);
   U2468 : MUX2_X1 port map( A => REGISTERS_18_13_port, B => n2830, S => n12, Z
                           => n1572);
   U2469 : MUX2_X1 port map( A => REGISTERS_18_12_port, B => n2831, S => n12, Z
                           => n1571);
   U2470 : MUX2_X1 port map( A => REGISTERS_18_11_port, B => n2832, S => n12, Z
                           => n1570);
   U2471 : MUX2_X1 port map( A => REGISTERS_18_10_port, B => n2833, S => n12, Z
                           => n1569);
   U2472 : MUX2_X1 port map( A => REGISTERS_18_9_port, B => n2834, S => n12, Z 
                           => n1568);
   U2473 : MUX2_X1 port map( A => REGISTERS_18_8_port, B => n2835, S => n12, Z 
                           => n1567);
   U2474 : MUX2_X1 port map( A => REGISTERS_18_7_port, B => n2836, S => n12, Z 
                           => n1566);
   U2475 : MUX2_X1 port map( A => REGISTERS_18_6_port, B => n2837, S => n12, Z 
                           => n1565);
   U2476 : MUX2_X1 port map( A => REGISTERS_18_5_port, B => n2838, S => n12, Z 
                           => n1564);
   U2477 : MUX2_X1 port map( A => REGISTERS_18_4_port, B => n2839, S => n12, Z 
                           => n1563);
   U2478 : MUX2_X1 port map( A => REGISTERS_18_3_port, B => n2840, S => n12, Z 
                           => n1562);
   U2479 : MUX2_X1 port map( A => REGISTERS_18_2_port, B => n2841, S => n12, Z 
                           => n1561);
   U2480 : MUX2_X1 port map( A => REGISTERS_18_1_port, B => n2842, S => n12, Z 
                           => n1560);
   U2481 : MUX2_X1 port map( A => REGISTERS_18_0_port, B => n2843, S => n12, Z 
                           => n1559);
   U2482 : OAI21_X1 port map( B1 => n2849, B2 => n2873, A => n274, ZN => n2875)
                           ;
   U2483 : MUX2_X1 port map( A => REGISTERS_19_31_port, B => n2811, S => n14, Z
                           => n1558);
   U2484 : MUX2_X1 port map( A => REGISTERS_19_30_port, B => n2813, S => n14, Z
                           => n1557);
   U2485 : MUX2_X1 port map( A => REGISTERS_19_29_port, B => n2814, S => n14, Z
                           => n1556);
   U2486 : MUX2_X1 port map( A => REGISTERS_19_28_port, B => n2815, S => n14, Z
                           => n1555);
   U2487 : MUX2_X1 port map( A => REGISTERS_19_27_port, B => n2816, S => n14, Z
                           => n1554);
   U2488 : MUX2_X1 port map( A => REGISTERS_19_26_port, B => n2817, S => n14, Z
                           => n1553);
   U2489 : MUX2_X1 port map( A => REGISTERS_19_25_port, B => n2818, S => n14, Z
                           => n1552);
   U2490 : MUX2_X1 port map( A => REGISTERS_19_24_port, B => n2819, S => n14, Z
                           => n1551);
   U2491 : MUX2_X1 port map( A => REGISTERS_19_23_port, B => n2820, S => n14, Z
                           => n1550);
   U2492 : MUX2_X1 port map( A => REGISTERS_19_22_port, B => n2821, S => n14, Z
                           => n1549);
   U2493 : MUX2_X1 port map( A => REGISTERS_19_21_port, B => n2822, S => n14, Z
                           => n1548);
   U2494 : MUX2_X1 port map( A => REGISTERS_19_20_port, B => n2823, S => n14, Z
                           => n1547);
   U2495 : MUX2_X1 port map( A => REGISTERS_19_19_port, B => n2824, S => n14, Z
                           => n1546);
   U2496 : MUX2_X1 port map( A => REGISTERS_19_18_port, B => n2825, S => n14, Z
                           => n1545);
   U2497 : MUX2_X1 port map( A => REGISTERS_19_17_port, B => n2826, S => n14, Z
                           => n1544);
   U2498 : MUX2_X1 port map( A => REGISTERS_19_16_port, B => n2827, S => n14, Z
                           => n1543);
   U2499 : MUX2_X1 port map( A => REGISTERS_19_15_port, B => n2828, S => n14, Z
                           => n1542);
   U2500 : MUX2_X1 port map( A => REGISTERS_19_14_port, B => n2829, S => n14, Z
                           => n1541);
   U2501 : MUX2_X1 port map( A => REGISTERS_19_13_port, B => n2830, S => n14, Z
                           => n1540);
   U2502 : MUX2_X1 port map( A => REGISTERS_19_12_port, B => n2831, S => n14, Z
                           => n1539);
   U2503 : MUX2_X1 port map( A => REGISTERS_19_11_port, B => n2832, S => n14, Z
                           => n1538);
   U2504 : MUX2_X1 port map( A => REGISTERS_19_10_port, B => n2833, S => n14, Z
                           => n1537);
   U2505 : MUX2_X1 port map( A => REGISTERS_19_9_port, B => n2834, S => n14, Z 
                           => n1536);
   U2506 : MUX2_X1 port map( A => REGISTERS_19_8_port, B => n2835, S => n14, Z 
                           => n1535);
   U2507 : MUX2_X1 port map( A => REGISTERS_19_7_port, B => n2836, S => n14, Z 
                           => n1534);
   U2508 : MUX2_X1 port map( A => REGISTERS_19_6_port, B => n2837, S => n14, Z 
                           => n1533);
   U2509 : MUX2_X1 port map( A => REGISTERS_19_5_port, B => n2838, S => n14, Z 
                           => n1532);
   U2510 : MUX2_X1 port map( A => REGISTERS_19_4_port, B => n2839, S => n14, Z 
                           => n1531);
   U2511 : MUX2_X1 port map( A => REGISTERS_19_3_port, B => n2840, S => n14, Z 
                           => n1530);
   U2512 : MUX2_X1 port map( A => REGISTERS_19_2_port, B => n2841, S => n14, Z 
                           => n1529);
   U2513 : MUX2_X1 port map( A => REGISTERS_19_1_port, B => n2842, S => n14, Z 
                           => n1528);
   U2514 : MUX2_X1 port map( A => REGISTERS_19_0_port, B => n2843, S => n14, Z 
                           => n1527);
   U2515 : OAI21_X1 port map( B1 => n2851, B2 => n2873, A => n274, ZN => n2876)
                           ;
   U2516 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => n2811, S => n16, Z
                           => n1526);
   U2517 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => n2813, S => n16, Z
                           => n1525);
   U2518 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => n2814, S => n16, Z
                           => n1524);
   U2519 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => n2815, S => n16, Z
                           => n1523);
   U2520 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => n2816, S => n16, Z
                           => n1522);
   U2521 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => n2817, S => n16, Z
                           => n1521);
   U2522 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => n2818, S => n16, Z
                           => n1520);
   U2523 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => n2819, S => n16, Z
                           => n1519);
   U2524 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => n2820, S => n16, Z
                           => n1518);
   U2525 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => n2821, S => n16, Z
                           => n1517);
   U2526 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => n2822, S => n16, Z
                           => n1516);
   U2527 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => n2823, S => n16, Z
                           => n1515);
   U2528 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => n2824, S => n16, Z
                           => n1514);
   U2529 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => n2825, S => n16, Z
                           => n1513);
   U2530 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => n2826, S => n16, Z
                           => n1512);
   U2531 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => n2827, S => n16, Z
                           => n1511);
   U2532 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => n2828, S => n16, Z
                           => n1510);
   U2533 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => n2829, S => n16, Z
                           => n1509);
   U2534 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => n2830, S => n16, Z
                           => n1508);
   U2535 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => n2831, S => n16, Z
                           => n1507);
   U2536 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => n2832, S => n16, Z
                           => n1506);
   U2537 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => n2833, S => n16, Z
                           => n1505);
   U2538 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => n2834, S => n16, Z 
                           => n1504);
   U2539 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => n2835, S => n16, Z 
                           => n1503);
   U2540 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => n2836, S => n16, Z 
                           => n1502);
   U2541 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => n2837, S => n16, Z 
                           => n1501);
   U2542 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => n2838, S => n16, Z 
                           => n1500);
   U2543 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => n2839, S => n16, Z 
                           => n1499);
   U2544 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => n2840, S => n16, Z 
                           => n1498);
   U2545 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => n2841, S => n16, Z 
                           => n1497);
   U2546 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => n2842, S => n16, Z 
                           => n1496);
   U2547 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => n2843, S => n16, Z 
                           => n1495);
   U2548 : OAI21_X1 port map( B1 => n2853, B2 => n2873, A => n274, ZN => n2877)
                           ;
   U2549 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => n2811, S => n18, Z
                           => n1494);
   U2550 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => n2813, S => n18, Z
                           => n1493);
   U2551 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => n2814, S => n18, Z
                           => n1492);
   U2552 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => n2815, S => n18, Z
                           => n1491);
   U2553 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => n2816, S => n18, Z
                           => n1490);
   U2554 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => n2817, S => n18, Z
                           => n1489);
   U2555 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => n2818, S => n18, Z
                           => n1488);
   U2556 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => n2819, S => n18, Z
                           => n1487);
   U2557 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => n2820, S => n18, Z
                           => n1486);
   U2558 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => n2821, S => n18, Z
                           => n1485);
   U2559 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => n2822, S => n18, Z
                           => n1484);
   U2560 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => n2823, S => n18, Z
                           => n1483);
   U2561 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => n2824, S => n18, Z
                           => n1482);
   U2562 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => n2825, S => n18, Z
                           => n1481);
   U2563 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => n2826, S => n18, Z
                           => n1480);
   U2564 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => n2827, S => n18, Z
                           => n1479);
   U2565 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => n2828, S => n18, Z
                           => n1478);
   U2566 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => n2829, S => n18, Z
                           => n1477);
   U2567 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => n2830, S => n18, Z
                           => n1476);
   U2568 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => n2831, S => n18, Z
                           => n1475);
   U2569 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => n2832, S => n18, Z
                           => n1474);
   U2570 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => n2833, S => n18, Z
                           => n1473);
   U2571 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => n2834, S => n18, Z 
                           => n1472);
   U2572 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => n2835, S => n18, Z 
                           => n1471);
   U2573 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => n2836, S => n18, Z 
                           => n1470);
   U2574 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => n2837, S => n18, Z 
                           => n1469);
   U2575 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => n2838, S => n18, Z 
                           => n1468);
   U2576 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => n2839, S => n18, Z 
                           => n1467);
   U2577 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => n2840, S => n18, Z 
                           => n1466);
   U2578 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => n2841, S => n18, Z 
                           => n1465);
   U2579 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => n2842, S => n18, Z 
                           => n1464);
   U2580 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => n2843, S => n18, Z 
                           => n1463);
   U2581 : OAI21_X1 port map( B1 => n2855, B2 => n2873, A => n274, ZN => n2878)
                           ;
   U2582 : MUX2_X1 port map( A => REGISTERS_22_31_port, B => n2811, S => n20, Z
                           => n1462);
   U2583 : MUX2_X1 port map( A => REGISTERS_22_30_port, B => n2813, S => n20, Z
                           => n1461);
   U2584 : MUX2_X1 port map( A => REGISTERS_22_29_port, B => n2814, S => n20, Z
                           => n1460);
   U2585 : MUX2_X1 port map( A => REGISTERS_22_28_port, B => n2815, S => n20, Z
                           => n1459);
   U2586 : MUX2_X1 port map( A => REGISTERS_22_27_port, B => n2816, S => n20, Z
                           => n1458);
   U2587 : MUX2_X1 port map( A => REGISTERS_22_26_port, B => n2817, S => n20, Z
                           => n1457);
   U2588 : MUX2_X1 port map( A => REGISTERS_22_25_port, B => n2818, S => n20, Z
                           => n1456);
   U2589 : MUX2_X1 port map( A => REGISTERS_22_24_port, B => n2819, S => n20, Z
                           => n1455);
   U2590 : MUX2_X1 port map( A => REGISTERS_22_23_port, B => n2820, S => n20, Z
                           => n1454);
   U2591 : MUX2_X1 port map( A => REGISTERS_22_22_port, B => n2821, S => n20, Z
                           => n1453);
   U2592 : MUX2_X1 port map( A => REGISTERS_22_21_port, B => n2822, S => n20, Z
                           => n1452);
   U2593 : MUX2_X1 port map( A => REGISTERS_22_20_port, B => n2823, S => n20, Z
                           => n1451);
   U2594 : MUX2_X1 port map( A => REGISTERS_22_19_port, B => n2824, S => n20, Z
                           => n1450);
   U2595 : MUX2_X1 port map( A => REGISTERS_22_18_port, B => n2825, S => n20, Z
                           => n1449);
   U2596 : MUX2_X1 port map( A => REGISTERS_22_17_port, B => n2826, S => n20, Z
                           => n1448);
   U2597 : MUX2_X1 port map( A => REGISTERS_22_16_port, B => n2827, S => n20, Z
                           => n1447);
   U2598 : MUX2_X1 port map( A => REGISTERS_22_15_port, B => n2828, S => n20, Z
                           => n1446);
   U2599 : MUX2_X1 port map( A => REGISTERS_22_14_port, B => n2829, S => n20, Z
                           => n1445);
   U2600 : MUX2_X1 port map( A => REGISTERS_22_13_port, B => n2830, S => n20, Z
                           => n1444);
   U2601 : MUX2_X1 port map( A => REGISTERS_22_12_port, B => n2831, S => n20, Z
                           => n1443);
   U2602 : MUX2_X1 port map( A => REGISTERS_22_11_port, B => n2832, S => n20, Z
                           => n1442);
   U2603 : MUX2_X1 port map( A => REGISTERS_22_10_port, B => n2833, S => n20, Z
                           => n1441);
   U2604 : MUX2_X1 port map( A => REGISTERS_22_9_port, B => n2834, S => n20, Z 
                           => n1440);
   U2605 : MUX2_X1 port map( A => REGISTERS_22_8_port, B => n2835, S => n20, Z 
                           => n1439);
   U2606 : MUX2_X1 port map( A => REGISTERS_22_7_port, B => n2836, S => n20, Z 
                           => n1438);
   U2607 : MUX2_X1 port map( A => REGISTERS_22_6_port, B => n2837, S => n20, Z 
                           => n1437);
   U2608 : MUX2_X1 port map( A => REGISTERS_22_5_port, B => n2838, S => n20, Z 
                           => n1436);
   U2609 : MUX2_X1 port map( A => REGISTERS_22_4_port, B => n2839, S => n20, Z 
                           => n1435);
   U2610 : MUX2_X1 port map( A => REGISTERS_22_3_port, B => n2840, S => n20, Z 
                           => n1434);
   U2611 : MUX2_X1 port map( A => REGISTERS_22_2_port, B => n2841, S => n20, Z 
                           => n1433);
   U2612 : MUX2_X1 port map( A => REGISTERS_22_1_port, B => n2842, S => n20, Z 
                           => n1432);
   U2613 : MUX2_X1 port map( A => REGISTERS_22_0_port, B => n2843, S => n20, Z 
                           => n1431);
   U2614 : OAI21_X1 port map( B1 => n2857, B2 => n2873, A => n274, ZN => n2879)
                           ;
   U2615 : MUX2_X1 port map( A => REGISTERS_23_31_port, B => n2811, S => n22, Z
                           => n1430);
   U2616 : MUX2_X1 port map( A => REGISTERS_23_30_port, B => n2813, S => n22, Z
                           => n1429);
   U2617 : MUX2_X1 port map( A => REGISTERS_23_29_port, B => n2814, S => n22, Z
                           => n1428);
   U2618 : MUX2_X1 port map( A => REGISTERS_23_28_port, B => n2815, S => n22, Z
                           => n1427);
   U2619 : MUX2_X1 port map( A => REGISTERS_23_27_port, B => n2816, S => n22, Z
                           => n1426);
   U2620 : MUX2_X1 port map( A => REGISTERS_23_26_port, B => n2817, S => n22, Z
                           => n1425);
   U2621 : MUX2_X1 port map( A => REGISTERS_23_25_port, B => n2818, S => n22, Z
                           => n1424);
   U2622 : MUX2_X1 port map( A => REGISTERS_23_24_port, B => n2819, S => n22, Z
                           => n1423);
   U2623 : MUX2_X1 port map( A => REGISTERS_23_23_port, B => n2820, S => n22, Z
                           => n1422);
   U2624 : MUX2_X1 port map( A => REGISTERS_23_22_port, B => n2821, S => n22, Z
                           => n1421);
   U2625 : MUX2_X1 port map( A => REGISTERS_23_21_port, B => n2822, S => n22, Z
                           => n1420);
   U2626 : MUX2_X1 port map( A => REGISTERS_23_20_port, B => n2823, S => n22, Z
                           => n1419);
   U2627 : MUX2_X1 port map( A => REGISTERS_23_19_port, B => n2824, S => n22, Z
                           => n1418);
   U2628 : MUX2_X1 port map( A => REGISTERS_23_18_port, B => n2825, S => n22, Z
                           => n1417);
   U2629 : MUX2_X1 port map( A => REGISTERS_23_17_port, B => n2826, S => n22, Z
                           => n1416);
   U2630 : MUX2_X1 port map( A => REGISTERS_23_16_port, B => n2827, S => n22, Z
                           => n1415);
   U2631 : MUX2_X1 port map( A => REGISTERS_23_15_port, B => n2828, S => n22, Z
                           => n1414);
   U2632 : MUX2_X1 port map( A => REGISTERS_23_14_port, B => n2829, S => n22, Z
                           => n1413);
   U2633 : MUX2_X1 port map( A => REGISTERS_23_13_port, B => n2830, S => n22, Z
                           => n1412);
   U2634 : MUX2_X1 port map( A => REGISTERS_23_12_port, B => n2831, S => n22, Z
                           => n1411);
   U2635 : MUX2_X1 port map( A => REGISTERS_23_11_port, B => n2832, S => n22, Z
                           => n1410);
   U2636 : MUX2_X1 port map( A => REGISTERS_23_10_port, B => n2833, S => n22, Z
                           => n1409);
   U2637 : MUX2_X1 port map( A => REGISTERS_23_9_port, B => n2834, S => n22, Z 
                           => n1408);
   U2638 : MUX2_X1 port map( A => REGISTERS_23_8_port, B => n2835, S => n22, Z 
                           => n1407);
   U2639 : MUX2_X1 port map( A => REGISTERS_23_7_port, B => n2836, S => n22, Z 
                           => n1406);
   U2640 : MUX2_X1 port map( A => REGISTERS_23_6_port, B => n2837, S => n22, Z 
                           => n1405);
   U2641 : MUX2_X1 port map( A => REGISTERS_23_5_port, B => n2838, S => n22, Z 
                           => n1404);
   U2642 : MUX2_X1 port map( A => REGISTERS_23_4_port, B => n2839, S => n22, Z 
                           => n1403);
   U2643 : MUX2_X1 port map( A => REGISTERS_23_3_port, B => n2840, S => n22, Z 
                           => n1402);
   U2644 : MUX2_X1 port map( A => REGISTERS_23_2_port, B => n2841, S => n22, Z 
                           => n1401);
   U2645 : MUX2_X1 port map( A => REGISTERS_23_1_port, B => n2842, S => n22, Z 
                           => n1400);
   U2646 : MUX2_X1 port map( A => REGISTERS_23_0_port, B => n2843, S => n22, Z 
                           => n1399);
   U2647 : OAI21_X1 port map( B1 => n2859, B2 => n2873, A => n275, ZN => n2880)
                           ;
   U2648 : NAND3_X1 port map( A1 => n2862, A2 => n2860, A3 => ADD_WR(4), ZN => 
                           n2873);
   U2649 : INV_X1 port map( A => ADD_WR(3), ZN => n2860);
   U2650 : MUX2_X1 port map( A => REGISTERS_24_31_port, B => n2811, S => n24, Z
                           => n1398);
   U2651 : MUX2_X1 port map( A => REGISTERS_24_30_port, B => n2813, S => n24, Z
                           => n1397);
   U2652 : MUX2_X1 port map( A => REGISTERS_24_29_port, B => n2814, S => n24, Z
                           => n1396);
   U2653 : MUX2_X1 port map( A => REGISTERS_24_28_port, B => n2815, S => n24, Z
                           => n1395);
   U2654 : MUX2_X1 port map( A => REGISTERS_24_27_port, B => n2816, S => n24, Z
                           => n1394);
   U2655 : MUX2_X1 port map( A => REGISTERS_24_26_port, B => n2817, S => n24, Z
                           => n1393);
   U2656 : MUX2_X1 port map( A => REGISTERS_24_25_port, B => n2818, S => n24, Z
                           => n1392);
   U2657 : MUX2_X1 port map( A => REGISTERS_24_24_port, B => n2819, S => n24, Z
                           => n1391);
   U2658 : MUX2_X1 port map( A => REGISTERS_24_23_port, B => n2820, S => n24, Z
                           => n1390);
   U2659 : MUX2_X1 port map( A => REGISTERS_24_22_port, B => n2821, S => n24, Z
                           => n1389);
   U2660 : MUX2_X1 port map( A => REGISTERS_24_21_port, B => n2822, S => n24, Z
                           => n1388);
   U2661 : MUX2_X1 port map( A => REGISTERS_24_20_port, B => n2823, S => n24, Z
                           => n1387);
   U2662 : MUX2_X1 port map( A => REGISTERS_24_19_port, B => n2824, S => n24, Z
                           => n1386);
   U2663 : MUX2_X1 port map( A => REGISTERS_24_18_port, B => n2825, S => n24, Z
                           => n1385);
   U2664 : MUX2_X1 port map( A => REGISTERS_24_17_port, B => n2826, S => n24, Z
                           => n1384);
   U2665 : MUX2_X1 port map( A => REGISTERS_24_16_port, B => n2827, S => n24, Z
                           => n1383);
   U2666 : MUX2_X1 port map( A => REGISTERS_24_15_port, B => n2828, S => n24, Z
                           => n1382);
   U2667 : MUX2_X1 port map( A => REGISTERS_24_14_port, B => n2829, S => n24, Z
                           => n1381);
   U2668 : MUX2_X1 port map( A => REGISTERS_24_13_port, B => n2830, S => n24, Z
                           => n1380);
   U2669 : MUX2_X1 port map( A => REGISTERS_24_12_port, B => n2831, S => n24, Z
                           => n1379);
   U2670 : MUX2_X1 port map( A => REGISTERS_24_11_port, B => n2832, S => n24, Z
                           => n1378);
   U2671 : MUX2_X1 port map( A => REGISTERS_24_10_port, B => n2833, S => n24, Z
                           => n1377);
   U2672 : MUX2_X1 port map( A => REGISTERS_24_9_port, B => n2834, S => n24, Z 
                           => n1376);
   U2673 : MUX2_X1 port map( A => REGISTERS_24_8_port, B => n2835, S => n24, Z 
                           => n1375);
   U2674 : MUX2_X1 port map( A => REGISTERS_24_7_port, B => n2836, S => n24, Z 
                           => n1374);
   U2675 : MUX2_X1 port map( A => REGISTERS_24_6_port, B => n2837, S => n24, Z 
                           => n1373);
   U2676 : MUX2_X1 port map( A => REGISTERS_24_5_port, B => n2838, S => n24, Z 
                           => n1372);
   U2677 : MUX2_X1 port map( A => REGISTERS_24_4_port, B => n2839, S => n24, Z 
                           => n1371);
   U2678 : MUX2_X1 port map( A => REGISTERS_24_3_port, B => n2840, S => n24, Z 
                           => n1370);
   U2679 : MUX2_X1 port map( A => REGISTERS_24_2_port, B => n2841, S => n24, Z 
                           => n1369);
   U2680 : MUX2_X1 port map( A => REGISTERS_24_1_port, B => n2842, S => n24, Z 
                           => n1368);
   U2681 : MUX2_X1 port map( A => REGISTERS_24_0_port, B => n2843, S => n24, Z 
                           => n1367);
   U2682 : OAI21_X1 port map( B1 => n2845, B2 => n2882, A => n275, ZN => n2881)
                           ;
   U2683 : NAND3_X1 port map( A1 => n2883, A2 => n2884, A3 => n2885, ZN => 
                           n2845);
   U2684 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => n2811, S => n26, Z
                           => n1366);
   U2685 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => n2813, S => n26, Z
                           => n1365);
   U2686 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => n2814, S => n26, Z
                           => n1364);
   U2687 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => n2815, S => n26, Z
                           => n1363);
   U2688 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => n2816, S => n26, Z
                           => n1362);
   U2689 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => n2817, S => n26, Z
                           => n1361);
   U2690 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => n2818, S => n26, Z
                           => n1360);
   U2691 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => n2819, S => n26, Z
                           => n1359);
   U2692 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => n2820, S => n26, Z
                           => n1358);
   U2693 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => n2821, S => n26, Z
                           => n1357);
   U2694 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => n2822, S => n26, Z
                           => n1356);
   U2695 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => n2823, S => n26, Z
                           => n1355);
   U2696 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => n2824, S => n26, Z
                           => n1354);
   U2697 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => n2825, S => n26, Z
                           => n1353);
   U2698 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => n2826, S => n26, Z
                           => n1352);
   U2699 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => n2827, S => n26, Z
                           => n1351);
   U2700 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => n2828, S => n26, Z
                           => n1350);
   U2701 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => n2829, S => n26, Z
                           => n1349);
   U2702 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => n2830, S => n26, Z
                           => n1348);
   U2703 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => n2831, S => n26, Z
                           => n1347);
   U2704 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => n2832, S => n26, Z
                           => n1346);
   U2705 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => n2833, S => n26, Z
                           => n1345);
   U2706 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => n2834, S => n26, Z 
                           => n1344);
   U2707 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => n2835, S => n26, Z 
                           => n1343);
   U2708 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => n2836, S => n26, Z 
                           => n1342);
   U2709 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => n2837, S => n26, Z 
                           => n1341);
   U2710 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => n2838, S => n26, Z 
                           => n1340);
   U2711 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => n2839, S => n26, Z 
                           => n1339);
   U2712 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => n2840, S => n26, Z 
                           => n1338);
   U2713 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => n2841, S => n26, Z 
                           => n1337);
   U2714 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => n2842, S => n26, Z 
                           => n1336);
   U2715 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => n2843, S => n26, Z 
                           => n1335);
   U2716 : OAI21_X1 port map( B1 => n2847, B2 => n2882, A => n275, ZN => n2886)
                           ;
   U2717 : NAND3_X1 port map( A1 => n2883, A2 => n2884, A3 => ADD_WR(0), ZN => 
                           n2847);
   U2718 : MUX2_X1 port map( A => REGISTERS_26_31_port, B => n2811, S => n28, Z
                           => n1334);
   U2719 : MUX2_X1 port map( A => REGISTERS_26_30_port, B => n2813, S => n28, Z
                           => n1333);
   U2720 : MUX2_X1 port map( A => REGISTERS_26_29_port, B => n2814, S => n28, Z
                           => n1332);
   U2721 : MUX2_X1 port map( A => REGISTERS_26_28_port, B => n2815, S => n28, Z
                           => n1331);
   U2722 : MUX2_X1 port map( A => REGISTERS_26_27_port, B => n2816, S => n28, Z
                           => n1330);
   U2723 : MUX2_X1 port map( A => REGISTERS_26_26_port, B => n2817, S => n28, Z
                           => n1329);
   U2724 : MUX2_X1 port map( A => REGISTERS_26_25_port, B => n2818, S => n28, Z
                           => n1328);
   U2725 : MUX2_X1 port map( A => REGISTERS_26_24_port, B => n2819, S => n28, Z
                           => n1327);
   U2726 : MUX2_X1 port map( A => REGISTERS_26_23_port, B => n2820, S => n28, Z
                           => n1326);
   U2727 : MUX2_X1 port map( A => REGISTERS_26_22_port, B => n2821, S => n28, Z
                           => n1325);
   U2728 : MUX2_X1 port map( A => REGISTERS_26_21_port, B => n2822, S => n28, Z
                           => n1324);
   U2729 : MUX2_X1 port map( A => REGISTERS_26_20_port, B => n2823, S => n28, Z
                           => n1323);
   U2730 : MUX2_X1 port map( A => REGISTERS_26_19_port, B => n2824, S => n28, Z
                           => n1322);
   U2731 : MUX2_X1 port map( A => REGISTERS_26_18_port, B => n2825, S => n28, Z
                           => n1321);
   U2732 : MUX2_X1 port map( A => REGISTERS_26_17_port, B => n2826, S => n28, Z
                           => n1320);
   U2733 : MUX2_X1 port map( A => REGISTERS_26_16_port, B => n2827, S => n28, Z
                           => n1319);
   U2734 : MUX2_X1 port map( A => REGISTERS_26_15_port, B => n2828, S => n28, Z
                           => n1318);
   U2735 : MUX2_X1 port map( A => REGISTERS_26_14_port, B => n2829, S => n28, Z
                           => n1317);
   U2736 : MUX2_X1 port map( A => REGISTERS_26_13_port, B => n2830, S => n28, Z
                           => n1316);
   U2737 : MUX2_X1 port map( A => REGISTERS_26_12_port, B => n2831, S => n28, Z
                           => n1315);
   U2738 : MUX2_X1 port map( A => REGISTERS_26_11_port, B => n2832, S => n28, Z
                           => n1314);
   U2739 : MUX2_X1 port map( A => REGISTERS_26_10_port, B => n2833, S => n28, Z
                           => n1313);
   U2740 : MUX2_X1 port map( A => REGISTERS_26_9_port, B => n2834, S => n28, Z 
                           => n1312);
   U2741 : MUX2_X1 port map( A => REGISTERS_26_8_port, B => n2835, S => n28, Z 
                           => n1311);
   U2742 : MUX2_X1 port map( A => REGISTERS_26_7_port, B => n2836, S => n28, Z 
                           => n1310);
   U2743 : MUX2_X1 port map( A => REGISTERS_26_6_port, B => n2837, S => n28, Z 
                           => n1309);
   U2744 : MUX2_X1 port map( A => REGISTERS_26_5_port, B => n2838, S => n28, Z 
                           => n1308);
   U2745 : MUX2_X1 port map( A => REGISTERS_26_4_port, B => n2839, S => n28, Z 
                           => n1307);
   U2746 : MUX2_X1 port map( A => REGISTERS_26_3_port, B => n2840, S => n28, Z 
                           => n1306);
   U2747 : MUX2_X1 port map( A => REGISTERS_26_2_port, B => n2841, S => n28, Z 
                           => n1305);
   U2748 : MUX2_X1 port map( A => REGISTERS_26_1_port, B => n2842, S => n28, Z 
                           => n1304);
   U2749 : MUX2_X1 port map( A => REGISTERS_26_0_port, B => n2843, S => n28, Z 
                           => n1303);
   U2750 : OAI21_X1 port map( B1 => n2849, B2 => n2882, A => n275, ZN => n2887)
                           ;
   U2751 : NAND3_X1 port map( A1 => n2885, A2 => n2884, A3 => ADD_WR(1), ZN => 
                           n2849);
   U2752 : MUX2_X1 port map( A => REGISTERS_27_31_port, B => n2811, S => n30, Z
                           => n1302);
   U2753 : MUX2_X1 port map( A => REGISTERS_27_30_port, B => n2813, S => n30, Z
                           => n1301);
   U2754 : MUX2_X1 port map( A => REGISTERS_27_29_port, B => n2814, S => n30, Z
                           => n1300);
   U2755 : MUX2_X1 port map( A => REGISTERS_27_28_port, B => n2815, S => n30, Z
                           => n1299);
   U2756 : MUX2_X1 port map( A => REGISTERS_27_27_port, B => n2816, S => n30, Z
                           => n1298);
   U2757 : MUX2_X1 port map( A => REGISTERS_27_26_port, B => n2817, S => n30, Z
                           => n1297);
   U2758 : MUX2_X1 port map( A => REGISTERS_27_25_port, B => n2818, S => n30, Z
                           => n1296);
   U2759 : MUX2_X1 port map( A => REGISTERS_27_24_port, B => n2819, S => n30, Z
                           => n1295);
   U2760 : MUX2_X1 port map( A => REGISTERS_27_23_port, B => n2820, S => n30, Z
                           => n1294);
   U2761 : MUX2_X1 port map( A => REGISTERS_27_22_port, B => n2821, S => n30, Z
                           => n1293);
   U2762 : MUX2_X1 port map( A => REGISTERS_27_21_port, B => n2822, S => n30, Z
                           => n1292);
   U2763 : MUX2_X1 port map( A => REGISTERS_27_20_port, B => n2823, S => n30, Z
                           => n1291);
   U2764 : MUX2_X1 port map( A => REGISTERS_27_19_port, B => n2824, S => n30, Z
                           => n1290);
   U2765 : MUX2_X1 port map( A => REGISTERS_27_18_port, B => n2825, S => n30, Z
                           => n1289);
   U2766 : MUX2_X1 port map( A => REGISTERS_27_17_port, B => n2826, S => n30, Z
                           => n1288);
   U2767 : MUX2_X1 port map( A => REGISTERS_27_16_port, B => n2827, S => n30, Z
                           => n1287);
   U2768 : MUX2_X1 port map( A => REGISTERS_27_15_port, B => n2828, S => n30, Z
                           => n1286);
   U2769 : MUX2_X1 port map( A => REGISTERS_27_14_port, B => n2829, S => n30, Z
                           => n1285);
   U2770 : MUX2_X1 port map( A => REGISTERS_27_13_port, B => n2830, S => n30, Z
                           => n1284);
   U2771 : MUX2_X1 port map( A => REGISTERS_27_12_port, B => n2831, S => n30, Z
                           => n1283);
   U2772 : MUX2_X1 port map( A => REGISTERS_27_11_port, B => n2832, S => n30, Z
                           => n1282);
   U2773 : MUX2_X1 port map( A => REGISTERS_27_10_port, B => n2833, S => n30, Z
                           => n1281);
   U2774 : MUX2_X1 port map( A => REGISTERS_27_9_port, B => n2834, S => n30, Z 
                           => n1280);
   U2775 : MUX2_X1 port map( A => REGISTERS_27_8_port, B => n2835, S => n30, Z 
                           => n1279);
   U2776 : MUX2_X1 port map( A => REGISTERS_27_7_port, B => n2836, S => n30, Z 
                           => n1278);
   U2777 : MUX2_X1 port map( A => REGISTERS_27_6_port, B => n2837, S => n30, Z 
                           => n1277);
   U2778 : MUX2_X1 port map( A => REGISTERS_27_5_port, B => n2838, S => n30, Z 
                           => n1276);
   U2779 : MUX2_X1 port map( A => REGISTERS_27_4_port, B => n2839, S => n30, Z 
                           => n1275);
   U2780 : MUX2_X1 port map( A => REGISTERS_27_3_port, B => n2840, S => n30, Z 
                           => n1274);
   U2781 : MUX2_X1 port map( A => REGISTERS_27_2_port, B => n2841, S => n30, Z 
                           => n1273);
   U2782 : MUX2_X1 port map( A => REGISTERS_27_1_port, B => n2842, S => n30, Z 
                           => n1272);
   U2783 : MUX2_X1 port map( A => REGISTERS_27_0_port, B => n2843, S => n30, Z 
                           => n1271);
   U2784 : OAI21_X1 port map( B1 => n2851, B2 => n2882, A => n275, ZN => n2888)
                           ;
   U2785 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2884, A3 => ADD_WR(1), ZN
                           => n2851);
   U2786 : INV_X1 port map( A => ADD_WR(2), ZN => n2884);
   U2787 : MUX2_X1 port map( A => REGISTERS_28_31_port, B => n2811, S => 
                           n32_port, Z => n1270);
   U2788 : MUX2_X1 port map( A => REGISTERS_28_30_port, B => n2813, S => 
                           n32_port, Z => n1269);
   U2789 : MUX2_X1 port map( A => REGISTERS_28_29_port, B => n2814, S => 
                           n32_port, Z => n1268);
   U2790 : MUX2_X1 port map( A => REGISTERS_28_28_port, B => n2815, S => 
                           n32_port, Z => n1267);
   U2791 : MUX2_X1 port map( A => REGISTERS_28_27_port, B => n2816, S => 
                           n32_port, Z => n1266);
   U2792 : MUX2_X1 port map( A => REGISTERS_28_26_port, B => n2817, S => 
                           n32_port, Z => n1265);
   U2793 : MUX2_X1 port map( A => REGISTERS_28_25_port, B => n2818, S => 
                           n32_port, Z => n1264);
   U2794 : MUX2_X1 port map( A => REGISTERS_28_24_port, B => n2819, S => 
                           n32_port, Z => n1263);
   U2795 : MUX2_X1 port map( A => REGISTERS_28_23_port, B => n2820, S => 
                           n32_port, Z => n1262);
   U2796 : MUX2_X1 port map( A => REGISTERS_28_22_port, B => n2821, S => 
                           n32_port, Z => n1261);
   U2797 : MUX2_X1 port map( A => REGISTERS_28_21_port, B => n2822, S => 
                           n32_port, Z => n1260);
   U2798 : MUX2_X1 port map( A => REGISTERS_28_20_port, B => n2823, S => 
                           n32_port, Z => n1259);
   U2799 : MUX2_X1 port map( A => REGISTERS_28_19_port, B => n2824, S => 
                           n32_port, Z => n1258);
   U2800 : MUX2_X1 port map( A => REGISTERS_28_18_port, B => n2825, S => 
                           n32_port, Z => n1257);
   U2801 : MUX2_X1 port map( A => REGISTERS_28_17_port, B => n2826, S => 
                           n32_port, Z => n1256);
   U2802 : MUX2_X1 port map( A => REGISTERS_28_16_port, B => n2827, S => 
                           n32_port, Z => n1255);
   U2803 : MUX2_X1 port map( A => REGISTERS_28_15_port, B => n2828, S => 
                           n32_port, Z => n1254);
   U2804 : MUX2_X1 port map( A => REGISTERS_28_14_port, B => n2829, S => 
                           n32_port, Z => n1253);
   U2805 : MUX2_X1 port map( A => REGISTERS_28_13_port, B => n2830, S => 
                           n32_port, Z => n1252);
   U2806 : MUX2_X1 port map( A => REGISTERS_28_12_port, B => n2831, S => 
                           n32_port, Z => n1251);
   U2807 : MUX2_X1 port map( A => REGISTERS_28_11_port, B => n2832, S => 
                           n32_port, Z => n1250);
   U2808 : MUX2_X1 port map( A => REGISTERS_28_10_port, B => n2833, S => 
                           n32_port, Z => n1249);
   U2809 : MUX2_X1 port map( A => REGISTERS_28_9_port, B => n2834, S => 
                           n32_port, Z => n1248);
   U2810 : MUX2_X1 port map( A => REGISTERS_28_8_port, B => n2835, S => 
                           n32_port, Z => n1247);
   U2811 : MUX2_X1 port map( A => REGISTERS_28_7_port, B => n2836, S => 
                           n32_port, Z => n1246);
   U2812 : MUX2_X1 port map( A => REGISTERS_28_6_port, B => n2837, S => 
                           n32_port, Z => n1245);
   U2813 : MUX2_X1 port map( A => REGISTERS_28_5_port, B => n2838, S => 
                           n32_port, Z => n1244);
   U2814 : MUX2_X1 port map( A => REGISTERS_28_4_port, B => n2839, S => 
                           n32_port, Z => n1243);
   U2815 : MUX2_X1 port map( A => REGISTERS_28_3_port, B => n2840, S => 
                           n32_port, Z => n1242);
   U2816 : MUX2_X1 port map( A => REGISTERS_28_2_port, B => n2841, S => 
                           n32_port, Z => n1241);
   U2817 : MUX2_X1 port map( A => REGISTERS_28_1_port, B => n2842, S => 
                           n32_port, Z => n1240);
   U2818 : MUX2_X1 port map( A => REGISTERS_28_0_port, B => n2843, S => 
                           n32_port, Z => n1239);
   U2819 : OAI21_X1 port map( B1 => n2853, B2 => n2882, A => n275, ZN => n2889)
                           ;
   U2820 : NAND3_X1 port map( A1 => n2885, A2 => n2883, A3 => ADD_WR(2), ZN => 
                           n2853);
   U2821 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => n2811, S => 
                           n34_port, Z => n1238);
   U2822 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => n2813, S => 
                           n34_port, Z => n1237);
   U2823 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => n2814, S => 
                           n34_port, Z => n1236);
   U2824 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => n2815, S => 
                           n34_port, Z => n1235);
   U2825 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => n2816, S => 
                           n34_port, Z => n1234);
   U2826 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => n2817, S => 
                           n34_port, Z => n1233);
   U2827 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => n2818, S => 
                           n34_port, Z => n1232);
   U2828 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => n2819, S => 
                           n34_port, Z => n1231);
   U2829 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => n2820, S => 
                           n34_port, Z => n1230);
   U2830 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => n2821, S => 
                           n34_port, Z => n1229);
   U2831 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => n2822, S => 
                           n34_port, Z => n1228);
   U2832 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => n2823, S => 
                           n34_port, Z => n1227);
   U2833 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => n2824, S => 
                           n34_port, Z => n1226);
   U2834 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => n2825, S => 
                           n34_port, Z => n1225);
   U2835 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => n2826, S => 
                           n34_port, Z => n1224);
   U2836 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => n2827, S => 
                           n34_port, Z => n1223);
   U2837 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => n2828, S => 
                           n34_port, Z => n1222);
   U2838 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => n2829, S => 
                           n34_port, Z => n1221);
   U2839 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => n2830, S => 
                           n34_port, Z => n1220);
   U2840 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => n2831, S => 
                           n34_port, Z => n1219);
   U2841 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => n2832, S => 
                           n34_port, Z => n1218);
   U2842 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => n2833, S => 
                           n34_port, Z => n1217);
   U2843 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => n2834, S => 
                           n34_port, Z => n1216);
   U2844 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => n2835, S => 
                           n34_port, Z => n1215);
   U2845 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => n2836, S => 
                           n34_port, Z => n1214);
   U2846 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => n2837, S => 
                           n34_port, Z => n1213);
   U2847 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => n2838, S => 
                           n34_port, Z => n1212);
   U2848 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => n2839, S => 
                           n34_port, Z => n1211);
   U2849 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => n2840, S => 
                           n34_port, Z => n1210);
   U2850 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => n2841, S => 
                           n34_port, Z => n1209);
   U2851 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => n2842, S => 
                           n34_port, Z => n1208);
   U2852 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => n2843, S => 
                           n34_port, Z => n1207);
   U2853 : OAI21_X1 port map( B1 => n2855, B2 => n2882, A => n275, ZN => n2890)
                           ;
   U2854 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2883, A3 => ADD_WR(2), ZN
                           => n2855);
   U2855 : INV_X1 port map( A => ADD_WR(1), ZN => n2883);
   U2856 : MUX2_X1 port map( A => REGISTERS_30_31_port, B => n2811, S => 
                           n36_port, Z => n1206);
   U2857 : MUX2_X1 port map( A => REGISTERS_30_30_port, B => n2813, S => 
                           n36_port, Z => n1205);
   U2858 : MUX2_X1 port map( A => REGISTERS_30_29_port, B => n2814, S => 
                           n36_port, Z => n1204);
   U2859 : MUX2_X1 port map( A => REGISTERS_30_28_port, B => n2815, S => 
                           n36_port, Z => n1203);
   U2860 : MUX2_X1 port map( A => REGISTERS_30_27_port, B => n2816, S => 
                           n36_port, Z => n1202);
   U2861 : MUX2_X1 port map( A => REGISTERS_30_26_port, B => n2817, S => 
                           n36_port, Z => n1201);
   U2862 : MUX2_X1 port map( A => REGISTERS_30_25_port, B => n2818, S => 
                           n36_port, Z => n1200);
   U2863 : MUX2_X1 port map( A => REGISTERS_30_24_port, B => n2819, S => 
                           n36_port, Z => n1199);
   U2864 : MUX2_X1 port map( A => REGISTERS_30_23_port, B => n2820, S => 
                           n36_port, Z => n1198);
   U2865 : MUX2_X1 port map( A => REGISTERS_30_22_port, B => n2821, S => 
                           n36_port, Z => n1197);
   U2866 : MUX2_X1 port map( A => REGISTERS_30_21_port, B => n2822, S => 
                           n36_port, Z => n1196);
   U2867 : MUX2_X1 port map( A => REGISTERS_30_20_port, B => n2823, S => 
                           n36_port, Z => n1195);
   U2868 : MUX2_X1 port map( A => REGISTERS_30_19_port, B => n2824, S => 
                           n36_port, Z => n1194);
   U2869 : MUX2_X1 port map( A => REGISTERS_30_18_port, B => n2825, S => 
                           n36_port, Z => n1193);
   U2870 : MUX2_X1 port map( A => REGISTERS_30_17_port, B => n2826, S => 
                           n36_port, Z => n1192);
   U2871 : MUX2_X1 port map( A => REGISTERS_30_16_port, B => n2827, S => 
                           n36_port, Z => n1191);
   U2872 : MUX2_X1 port map( A => REGISTERS_30_15_port, B => n2828, S => 
                           n36_port, Z => n1190);
   U2873 : MUX2_X1 port map( A => REGISTERS_30_14_port, B => n2829, S => 
                           n36_port, Z => n1189);
   U2874 : MUX2_X1 port map( A => REGISTERS_30_13_port, B => n2830, S => 
                           n36_port, Z => n1188);
   U2875 : MUX2_X1 port map( A => REGISTERS_30_12_port, B => n2831, S => 
                           n36_port, Z => n1187);
   U2876 : MUX2_X1 port map( A => REGISTERS_30_11_port, B => n2832, S => 
                           n36_port, Z => n1186);
   U2877 : MUX2_X1 port map( A => REGISTERS_30_10_port, B => n2833, S => 
                           n36_port, Z => n1185);
   U2878 : MUX2_X1 port map( A => REGISTERS_30_9_port, B => n2834, S => 
                           n36_port, Z => n1184);
   U2879 : MUX2_X1 port map( A => REGISTERS_30_8_port, B => n2835, S => 
                           n36_port, Z => n1183);
   U2880 : MUX2_X1 port map( A => REGISTERS_30_7_port, B => n2836, S => 
                           n36_port, Z => n1182);
   U2881 : MUX2_X1 port map( A => REGISTERS_30_6_port, B => n2837, S => 
                           n36_port, Z => n1181);
   U2882 : MUX2_X1 port map( A => REGISTERS_30_5_port, B => n2838, S => 
                           n36_port, Z => n1180);
   U2883 : MUX2_X1 port map( A => REGISTERS_30_4_port, B => n2839, S => 
                           n36_port, Z => n1179);
   U2884 : MUX2_X1 port map( A => REGISTERS_30_3_port, B => n2840, S => 
                           n36_port, Z => n1178);
   U2885 : MUX2_X1 port map( A => REGISTERS_30_2_port, B => n2841, S => 
                           n36_port, Z => n1177);
   U2886 : MUX2_X1 port map( A => REGISTERS_30_1_port, B => n2842, S => 
                           n36_port, Z => n1176);
   U2887 : MUX2_X1 port map( A => REGISTERS_30_0_port, B => n2843, S => 
                           n36_port, Z => n1175);
   U2888 : OAI21_X1 port map( B1 => n2857, B2 => n2882, A => n275, ZN => n2891)
                           ;
   U2889 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n2885, A3 => ADD_WR(2), ZN
                           => n2857);
   U2890 : INV_X1 port map( A => ADD_WR(0), ZN => n2885);
   U2891 : MUX2_X1 port map( A => REGISTERS_31_31_port, B => n2811, S => 
                           n38_port, Z => n1174);
   U2892 : AND2_X1 port map( A1 => DATAIN(31), A2 => n275, ZN => n2811);
   U2893 : MUX2_X1 port map( A => REGISTERS_31_30_port, B => n2813, S => 
                           n38_port, Z => n1173);
   U2894 : AND2_X1 port map( A1 => DATAIN(30), A2 => n275, ZN => n2813);
   U2895 : MUX2_X1 port map( A => REGISTERS_31_29_port, B => n2814, S => 
                           n38_port, Z => n1172);
   U2896 : AND2_X1 port map( A1 => DATAIN(29), A2 => n275, ZN => n2814);
   U2897 : MUX2_X1 port map( A => REGISTERS_31_28_port, B => n2815, S => 
                           n38_port, Z => n1171);
   U2898 : AND2_X1 port map( A1 => DATAIN(28), A2 => n275, ZN => n2815);
   U2899 : MUX2_X1 port map( A => REGISTERS_31_27_port, B => n2816, S => 
                           n38_port, Z => n1170);
   U2900 : AND2_X1 port map( A1 => DATAIN(27), A2 => n276, ZN => n2816);
   U2901 : MUX2_X1 port map( A => REGISTERS_31_26_port, B => n2817, S => 
                           n38_port, Z => n1169);
   U2902 : AND2_X1 port map( A1 => DATAIN(26), A2 => n276, ZN => n2817);
   U2903 : MUX2_X1 port map( A => REGISTERS_31_25_port, B => n2818, S => 
                           n38_port, Z => n1168);
   U2904 : AND2_X1 port map( A1 => DATAIN(25), A2 => n276, ZN => n2818);
   U2905 : MUX2_X1 port map( A => REGISTERS_31_24_port, B => n2819, S => 
                           n38_port, Z => n1167);
   U2906 : AND2_X1 port map( A1 => DATAIN(24), A2 => n276, ZN => n2819);
   U2907 : MUX2_X1 port map( A => REGISTERS_31_23_port, B => n2820, S => 
                           n38_port, Z => n1166);
   U2908 : AND2_X1 port map( A1 => DATAIN(23), A2 => n276, ZN => n2820);
   U2909 : MUX2_X1 port map( A => REGISTERS_31_22_port, B => n2821, S => 
                           n38_port, Z => n1165);
   U2910 : AND2_X1 port map( A1 => DATAIN(22), A2 => n276, ZN => n2821);
   U2911 : MUX2_X1 port map( A => REGISTERS_31_21_port, B => n2822, S => 
                           n38_port, Z => n1164);
   U2912 : AND2_X1 port map( A1 => DATAIN(21), A2 => n276, ZN => n2822);
   U2913 : MUX2_X1 port map( A => REGISTERS_31_20_port, B => n2823, S => 
                           n38_port, Z => n1163);
   U2914 : AND2_X1 port map( A1 => DATAIN(20), A2 => n276, ZN => n2823);
   U2915 : MUX2_X1 port map( A => REGISTERS_31_19_port, B => n2824, S => 
                           n38_port, Z => n1162);
   U2916 : AND2_X1 port map( A1 => DATAIN(19), A2 => n276, ZN => n2824);
   U2917 : MUX2_X1 port map( A => REGISTERS_31_18_port, B => n2825, S => 
                           n38_port, Z => n1161);
   U2918 : AND2_X1 port map( A1 => DATAIN(18), A2 => n276, ZN => n2825);
   U2919 : MUX2_X1 port map( A => REGISTERS_31_17_port, B => n2826, S => 
                           n38_port, Z => n1160);
   U2920 : AND2_X1 port map( A1 => DATAIN(17), A2 => n276, ZN => n2826);
   U2921 : MUX2_X1 port map( A => REGISTERS_31_16_port, B => n2827, S => 
                           n38_port, Z => n1159);
   U2922 : AND2_X1 port map( A1 => DATAIN(16), A2 => n276, ZN => n2827);
   U2923 : MUX2_X1 port map( A => REGISTERS_31_15_port, B => n2828, S => 
                           n38_port, Z => n1158);
   U2924 : AND2_X1 port map( A1 => DATAIN(15), A2 => n276, ZN => n2828);
   U2925 : MUX2_X1 port map( A => REGISTERS_31_14_port, B => n2829, S => 
                           n38_port, Z => n1157);
   U2926 : AND2_X1 port map( A1 => DATAIN(14), A2 => n276, ZN => n2829);
   U2927 : MUX2_X1 port map( A => REGISTERS_31_13_port, B => n2830, S => 
                           n38_port, Z => n1156);
   U2928 : AND2_X1 port map( A1 => DATAIN(13), A2 => n275, ZN => n2830);
   U2929 : MUX2_X1 port map( A => REGISTERS_31_12_port, B => n2831, S => 
                           n38_port, Z => n1155);
   U2930 : AND2_X1 port map( A1 => DATAIN(12), A2 => n276, ZN => n2831);
   U2931 : MUX2_X1 port map( A => REGISTERS_31_11_port, B => n2832, S => 
                           n38_port, Z => n1154);
   U2932 : AND2_X1 port map( A1 => DATAIN(11), A2 => n276, ZN => n2832);
   U2933 : MUX2_X1 port map( A => REGISTERS_31_10_port, B => n2833, S => 
                           n38_port, Z => n1153);
   U2934 : AND2_X1 port map( A1 => DATAIN(10), A2 => n277, ZN => n2833);
   U2935 : MUX2_X1 port map( A => REGISTERS_31_9_port, B => n2834, S => 
                           n38_port, Z => n1152);
   U2936 : AND2_X1 port map( A1 => DATAIN(9), A2 => n277, ZN => n2834);
   U2937 : MUX2_X1 port map( A => REGISTERS_31_8_port, B => n2835, S => 
                           n38_port, Z => n1151);
   U2938 : AND2_X1 port map( A1 => DATAIN(8), A2 => n277, ZN => n2835);
   U2939 : MUX2_X1 port map( A => REGISTERS_31_7_port, B => n2836, S => 
                           n38_port, Z => n1150);
   U2940 : AND2_X1 port map( A1 => DATAIN(7), A2 => n277, ZN => n2836);
   U2941 : MUX2_X1 port map( A => REGISTERS_31_6_port, B => n2837, S => 
                           n38_port, Z => n1149);
   U2942 : AND2_X1 port map( A1 => DATAIN(6), A2 => n277, ZN => n2837);
   U2943 : MUX2_X1 port map( A => REGISTERS_31_5_port, B => n2838, S => 
                           n38_port, Z => n1148);
   U2944 : AND2_X1 port map( A1 => DATAIN(5), A2 => n277, ZN => n2838);
   U2945 : MUX2_X1 port map( A => REGISTERS_31_4_port, B => n2839, S => 
                           n38_port, Z => n1147);
   U2946 : AND2_X1 port map( A1 => DATAIN(4), A2 => n277, ZN => n2839);
   U2947 : MUX2_X1 port map( A => REGISTERS_31_3_port, B => n2840, S => 
                           n38_port, Z => n1146);
   U2948 : AND2_X1 port map( A1 => DATAIN(3), A2 => n277, ZN => n2840);
   U2949 : MUX2_X1 port map( A => REGISTERS_31_2_port, B => n2841, S => 
                           n38_port, Z => n1145);
   U2950 : AND2_X1 port map( A1 => DATAIN(2), A2 => n277, ZN => n2841);
   U2951 : MUX2_X1 port map( A => REGISTERS_31_1_port, B => n2842, S => 
                           n38_port, Z => n1144);
   U2952 : AND2_X1 port map( A1 => DATAIN(1), A2 => n277, ZN => n2842);
   U2953 : MUX2_X1 port map( A => REGISTERS_31_0_port, B => n2843, S => 
                           n38_port, Z => n1143);
   U2954 : OAI21_X1 port map( B1 => n2859, B2 => n2882, A => n273, ZN => n2892)
                           ;
   U2955 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n2862, A3 => ADD_WR(4), ZN
                           => n2882);
   U2956 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n2862);
   U2957 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n2859);
   U2958 : AND2_X1 port map( A1 => DATAIN(0), A2 => n277, ZN => n2843);
   U2959 : AND2_X1 port map( A1 => N96, A2 => n2893, ZN => N448);
   U2960 : AND2_X1 port map( A1 => N97, A2 => n2893, ZN => N447);
   U2961 : AND2_X1 port map( A1 => N98, A2 => n2893, ZN => N446);
   U2962 : AND2_X1 port map( A1 => N99, A2 => n2893, ZN => N445);
   U2963 : AND2_X1 port map( A1 => N100, A2 => n2893, ZN => N444);
   U2964 : AND2_X1 port map( A1 => N101, A2 => n2893, ZN => N443);
   U2965 : AND2_X1 port map( A1 => N102, A2 => n2893, ZN => N442);
   U2966 : AND2_X1 port map( A1 => N103, A2 => n2893, ZN => N441);
   U2967 : AND2_X1 port map( A1 => N104, A2 => n2893, ZN => N440);
   U2968 : AND2_X1 port map( A1 => N105, A2 => n2893, ZN => N439);
   U2969 : AND2_X1 port map( A1 => N106, A2 => n2893, ZN => N438);
   U2970 : AND2_X1 port map( A1 => N107, A2 => n2893, ZN => N437);
   U2971 : AND2_X1 port map( A1 => N108, A2 => n2893, ZN => N436);
   U2972 : AND2_X1 port map( A1 => N109, A2 => n2893, ZN => N435);
   U2973 : AND2_X1 port map( A1 => N110, A2 => n2893, ZN => N434);
   U2974 : AND2_X1 port map( A1 => N111, A2 => n2893, ZN => N433);
   U2975 : AND2_X1 port map( A1 => N112, A2 => n2893, ZN => N432);
   U2976 : AND2_X1 port map( A1 => N113, A2 => n2893, ZN => N431);
   U2977 : AND2_X1 port map( A1 => N114, A2 => n2893, ZN => N430);
   U2978 : AND2_X1 port map( A1 => N115, A2 => n2893, ZN => N429);
   U2979 : AND2_X1 port map( A1 => N116, A2 => n2893, ZN => N428);
   U2980 : AND2_X1 port map( A1 => N117, A2 => n2893, ZN => N427);
   U2981 : AND2_X1 port map( A1 => N118, A2 => n2893, ZN => N426);
   U2982 : AND2_X1 port map( A1 => N119, A2 => n2893, ZN => N425);
   U2983 : AND2_X1 port map( A1 => N120, A2 => n2893, ZN => N424);
   U2984 : AND2_X1 port map( A1 => N121, A2 => n2893, ZN => N423);
   U2985 : AND2_X1 port map( A1 => N122, A2 => n2893, ZN => N422);
   U2986 : AND2_X1 port map( A1 => N123, A2 => n2893, ZN => N421);
   U2987 : AND2_X1 port map( A1 => N124, A2 => n2893, ZN => N420);
   U2988 : AND2_X1 port map( A1 => N125, A2 => n2893, ZN => N419);
   U2989 : AND2_X1 port map( A1 => N126, A2 => n2893, ZN => N418);
   U2990 : AND2_X1 port map( A1 => N127, A2 => n2893, ZN => N417);
   U2991 : AND3_X1 port map( A1 => ENABLE, A2 => n277, A3 => RD2, ZN => n2893);
   U2992 : AND2_X1 port map( A1 => N31, A2 => n2894, ZN => N416);
   U2993 : AND2_X1 port map( A1 => N32, A2 => n2894, ZN => N415);
   U2994 : AND2_X1 port map( A1 => N33, A2 => n2894, ZN => N414);
   U2995 : AND2_X1 port map( A1 => N34, A2 => n2894, ZN => N413);
   U2996 : AND2_X1 port map( A1 => N35, A2 => n2894, ZN => N412);
   U2997 : AND2_X1 port map( A1 => N36, A2 => n2894, ZN => N411);
   U2998 : AND2_X1 port map( A1 => N37, A2 => n2894, ZN => N410);
   U2999 : AND2_X1 port map( A1 => N38, A2 => n2894, ZN => N409);
   U3000 : AND2_X1 port map( A1 => N39, A2 => n2894, ZN => N408);
   U3001 : AND2_X1 port map( A1 => N40, A2 => n2894, ZN => N407);
   U3002 : AND2_X1 port map( A1 => N41, A2 => n2894, ZN => N406);
   U3003 : AND2_X1 port map( A1 => N42, A2 => n2894, ZN => N405);
   U3004 : AND2_X1 port map( A1 => N43, A2 => n2894, ZN => N404);
   U3005 : AND2_X1 port map( A1 => N44, A2 => n2894, ZN => N403);
   U3006 : AND2_X1 port map( A1 => N45, A2 => n2894, ZN => N402);
   U3007 : AND2_X1 port map( A1 => N46, A2 => n2894, ZN => N401);
   U3008 : AND2_X1 port map( A1 => N47, A2 => n2894, ZN => N400);
   U3009 : AND2_X1 port map( A1 => N48, A2 => n2894, ZN => N399);
   U3010 : AND2_X1 port map( A1 => N49, A2 => n2894, ZN => N398);
   U3011 : AND2_X1 port map( A1 => N50, A2 => n2894, ZN => N397);
   U3012 : AND2_X1 port map( A1 => N51, A2 => n2894, ZN => N396);
   U3013 : AND2_X1 port map( A1 => N52, A2 => n2894, ZN => N395);
   U3014 : AND2_X1 port map( A1 => N53, A2 => n2894, ZN => N394);
   U3015 : AND2_X1 port map( A1 => N54, A2 => n2894, ZN => N393);
   U3016 : AND2_X1 port map( A1 => N55, A2 => n2894, ZN => N392);
   U3017 : AND2_X1 port map( A1 => N56, A2 => n2894, ZN => N391);
   U3018 : AND2_X1 port map( A1 => N57, A2 => n2894, ZN => N390);
   U3019 : AND2_X1 port map( A1 => N58, A2 => n2894, ZN => N389);
   U3020 : AND2_X1 port map( A1 => N59, A2 => n2894, ZN => N388);
   U3021 : AND2_X1 port map( A1 => N60, A2 => n2894, ZN => N387);
   U3022 : AND2_X1 port map( A1 => N61, A2 => n2894, ZN => N386);
   U3023 : AND2_X1 port map( A1 => N62, A2 => n2894, ZN => N385);
   U3024 : AND3_X1 port map( A1 => ENABLE, A2 => n277, A3 => RD1, ZN => n2894);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n5_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  Q :
         out std_logic_vector (4 downto 0));

end reg_nbit_n5_0;

architecture SYN_struc of reg_nbit_n5_0 is

   component FD_2084
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2085
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2086
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2087
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2088
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;

begin
   
   D_I_0 : FD_2088 port map( D => d(0), CK => clk, RESET => reset, Q => Q(0));
   D_I_1 : FD_2087 port map( D => d(1), CK => clk, RESET => reset, Q => Q(1));
   D_I_2 : FD_2086 port map( D => d(2), CK => clk, RESET => reset, Q => Q(2));
   D_I_3 : FD_2085 port map( D => d(3), CK => clk, RESET => reset, Q => Q(3));
   D_I_4 : FD_2084 port map( D => d(4), CK => clk, RESET => reset, Q => Q(4));

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n32_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0);  Q 
         : out std_logic_vector (31 downto 0));

end reg_nbit_n32_0;

architecture SYN_struc of reg_nbit_n32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2153
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2154
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2155
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2156
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2157
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2158
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2159
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2160
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2161
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2162
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2163
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2164
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2165
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2166
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2167
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2168
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2169
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2170
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2171
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2172
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2173
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2174
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2175
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2176
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2177
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2178
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2179
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2180
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2181
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2182
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2183
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2184
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   D_I_0 : FD_2184 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_2183 port map( D => d(1), CK => n1, RESET => reset, Q => Q(1));
   D_I_2 : FD_2182 port map( D => d(2), CK => n1, RESET => reset, Q => Q(2));
   D_I_3 : FD_2181 port map( D => d(3), CK => n1, RESET => reset, Q => Q(3));
   D_I_4 : FD_2180 port map( D => d(4), CK => n1, RESET => reset, Q => Q(4));
   D_I_5 : FD_2179 port map( D => d(5), CK => n1, RESET => reset, Q => Q(5));
   D_I_6 : FD_2178 port map( D => d(6), CK => n1, RESET => reset, Q => Q(6));
   D_I_7 : FD_2177 port map( D => d(7), CK => n1, RESET => reset, Q => Q(7));
   D_I_8 : FD_2176 port map( D => d(8), CK => n1, RESET => reset, Q => Q(8));
   D_I_9 : FD_2175 port map( D => d(9), CK => n1, RESET => reset, Q => Q(9));
   D_I_10 : FD_2174 port map( D => d(10), CK => n1, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2173 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2172 port map( D => d(12), CK => n2, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2171 port map( D => d(13), CK => n2, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2170 port map( D => d(14), CK => n2, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2169 port map( D => d(15), CK => n2, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2168 port map( D => d(16), CK => n2, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2167 port map( D => d(17), CK => n2, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2166 port map( D => d(18), CK => n2, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2165 port map( D => d(19), CK => n2, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2164 port map( D => d(20), CK => n2, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2163 port map( D => d(21), CK => n2, RESET => reset, Q => Q(21))
                           ;
   D_I_22 : FD_2162 port map( D => d(22), CK => n3, RESET => reset, Q => Q(22))
                           ;
   D_I_23 : FD_2161 port map( D => d(23), CK => n3, RESET => reset, Q => Q(23))
                           ;
   D_I_24 : FD_2160 port map( D => d(24), CK => n3, RESET => reset, Q => Q(24))
                           ;
   D_I_25 : FD_2159 port map( D => d(25), CK => n3, RESET => reset, Q => Q(25))
                           ;
   D_I_26 : FD_2158 port map( D => d(26), CK => n3, RESET => reset, Q => Q(26))
                           ;
   D_I_27 : FD_2157 port map( D => d(27), CK => n3, RESET => reset, Q => Q(27))
                           ;
   D_I_28 : FD_2156 port map( D => d(28), CK => n3, RESET => reset, Q => Q(28))
                           ;
   D_I_29 : FD_2155 port map( D => d(29), CK => n3, RESET => reset, Q => Q(29))
                           ;
   D_I_30 : FD_2154 port map( D => d(30), CK => n3, RESET => reset, Q => Q(30))
                           ;
   D_I_31 : FD_2153 port map( D => d(31), CK => n3, RESET => reset, Q => Q(31))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n1);
   U2 : BUF_X1 port map( A => clk, Z => n2);
   U3 : BUF_X1 port map( A => clk, Z => n3);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FD_0 is

   port( D, CK, RESET : in std_logic;  Q : out std_logic);

end FD_0;

architecture SYN_PLUTO of FD_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n_5533 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => D, CK => CK, RN => n1, Q => Q, QN => n_5533);
   U3 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_PLUTO;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity write_back_stage_N32 is

   port( data_from_memory, data_from_alu : in std_logic_vector (31 downto 0);  
         data_to_rf : out std_logic_vector (31 downto 0);  select_wb : in 
         std_logic);

end write_back_stage_N32;

architecture SYN_structural of write_back_stage_N32 is

   component MUX_zbit_nbit_N32_Z1_1
      port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   wb_mux : MUX_zbit_nbit_N32_Z1_1 port map( inputs(0) => data_from_memory(31),
                           inputs(1) => data_from_memory(30), inputs(2) => 
                           data_from_memory(29), inputs(3) => 
                           data_from_memory(28), inputs(4) => 
                           data_from_memory(27), inputs(5) => 
                           data_from_memory(26), inputs(6) => 
                           data_from_memory(25), inputs(7) => 
                           data_from_memory(24), inputs(8) => 
                           data_from_memory(23), inputs(9) => 
                           data_from_memory(22), inputs(10) => 
                           data_from_memory(21), inputs(11) => 
                           data_from_memory(20), inputs(12) => 
                           data_from_memory(19), inputs(13) => 
                           data_from_memory(18), inputs(14) => 
                           data_from_memory(17), inputs(15) => 
                           data_from_memory(16), inputs(16) => 
                           data_from_memory(15), inputs(17) => 
                           data_from_memory(14), inputs(18) => 
                           data_from_memory(13), inputs(19) => 
                           data_from_memory(12), inputs(20) => 
                           data_from_memory(11), inputs(21) => 
                           data_from_memory(10), inputs(22) => 
                           data_from_memory(9), inputs(23) => 
                           data_from_memory(8), inputs(24) => 
                           data_from_memory(7), inputs(25) => 
                           data_from_memory(6), inputs(26) => 
                           data_from_memory(5), inputs(27) => 
                           data_from_memory(4), inputs(28) => 
                           data_from_memory(3), inputs(29) => 
                           data_from_memory(2), inputs(30) => 
                           data_from_memory(1), inputs(31) => 
                           data_from_memory(0), inputs(32) => data_from_alu(31)
                           , inputs(33) => data_from_alu(30), inputs(34) => 
                           data_from_alu(29), inputs(35) => data_from_alu(28), 
                           inputs(36) => data_from_alu(27), inputs(37) => 
                           data_from_alu(26), inputs(38) => data_from_alu(25), 
                           inputs(39) => data_from_alu(24), inputs(40) => 
                           data_from_alu(23), inputs(41) => data_from_alu(22), 
                           inputs(42) => data_from_alu(21), inputs(43) => 
                           data_from_alu(20), inputs(44) => data_from_alu(19), 
                           inputs(45) => data_from_alu(18), inputs(46) => 
                           data_from_alu(17), inputs(47) => data_from_alu(16), 
                           inputs(48) => data_from_alu(15), inputs(49) => 
                           data_from_alu(14), inputs(50) => data_from_alu(13), 
                           inputs(51) => data_from_alu(12), inputs(52) => 
                           data_from_alu(11), inputs(53) => data_from_alu(10), 
                           inputs(54) => data_from_alu(9), inputs(55) => 
                           data_from_alu(8), inputs(56) => data_from_alu(7), 
                           inputs(57) => data_from_alu(6), inputs(58) => 
                           data_from_alu(5), inputs(59) => data_from_alu(4), 
                           inputs(60) => data_from_alu(3), inputs(61) => 
                           data_from_alu(2), inputs(62) => data_from_alu(1), 
                           inputs(63) => data_from_alu(0), SEL => select_wb, 
                           Y(31) => data_to_rf(31), Y(30) => data_to_rf(30), 
                           Y(29) => data_to_rf(29), Y(28) => data_to_rf(28), 
                           Y(27) => data_to_rf(27), Y(26) => data_to_rf(26), 
                           Y(25) => data_to_rf(25), Y(24) => data_to_rf(24), 
                           Y(23) => data_to_rf(23), Y(22) => data_to_rf(22), 
                           Y(21) => data_to_rf(21), Y(20) => data_to_rf(20), 
                           Y(19) => data_to_rf(19), Y(18) => data_to_rf(18), 
                           Y(17) => data_to_rf(17), Y(16) => data_to_rf(16), 
                           Y(15) => data_to_rf(15), Y(14) => data_to_rf(14), 
                           Y(13) => data_to_rf(13), Y(12) => data_to_rf(12), 
                           Y(11) => data_to_rf(11), Y(10) => data_to_rf(10), 
                           Y(9) => data_to_rf(9), Y(8) => data_to_rf(8), Y(7) 
                           => data_to_rf(7), Y(6) => data_to_rf(6), Y(5) => 
                           data_to_rf(5), Y(4) => data_to_rf(4), Y(3) => 
                           data_to_rf(3), Y(2) => data_to_rf(2), Y(1) => 
                           data_to_rf(1), Y(0) => data_to_rf(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity memory_stage_N32_PC_SIZE32 is

   port( clk, rst : in std_logic;  new_pc_value : in std_logic_vector (31 
         downto 0);  new_pc_value_branch : out std_logic_vector (31 downto 0); 
         select_pc : in std_logic;  alu_output_val, value_to_mem : in 
         std_logic_vector (31 downto 0);  data_from_memory, data_from_alu : out
         std_logic_vector (31 downto 0);  dram_enable_cu, dram_r_nw_cu : in 
         std_logic;  dram_ready_cu : out std_logic;  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end memory_stage_N32_PC_SIZE32;

architecture SYN_structural of memory_stage_N32_PC_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component reg_nbit_n32_7
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_8
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX_zbit_nbit_N32_Z1_2
      port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, data_ir_31_port, data_ir_30_port, data_ir_29_port, 
      data_ir_28_port, data_ir_27_port, data_ir_26_port, data_ir_25_port, 
      data_ir_24_port, data_ir_23_port, data_ir_22_port, data_ir_21_port, 
      data_ir_20_port, data_ir_19_port, data_ir_18_port, data_ir_17_port, 
      data_ir_16_port, data_ir_15_port, data_ir_14_port, data_ir_13_port, 
      data_ir_12_port, data_ir_11_port, data_ir_10_port, data_ir_9_port, 
      data_ir_8_port, data_ir_7_port, data_ir_6_port, data_ir_5_port, 
      data_ir_4_port, data_ir_3_port, data_ir_2_port, data_ir_1_port, 
      data_ir_0_port, n2, n1, n3 : std_logic;

begin
   dram_ready_cu <= DRAM_READY;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, X_Logic0_port, X_Logic0_port );
   DRAM_ENABLE <= dram_enable_cu;
   DRAM_READNOTWRITE <= dram_r_nw_cu;
   
   X_Logic0_port <= '0';
   branch_mux : MUX_zbit_nbit_N32_Z1_2 port map( inputs(0) => new_pc_value(31),
                           inputs(1) => new_pc_value(30), inputs(2) => 
                           new_pc_value(29), inputs(3) => new_pc_value(28), 
                           inputs(4) => new_pc_value(27), inputs(5) => 
                           new_pc_value(26), inputs(6) => new_pc_value(25), 
                           inputs(7) => new_pc_value(24), inputs(8) => 
                           new_pc_value(23), inputs(9) => new_pc_value(22), 
                           inputs(10) => new_pc_value(21), inputs(11) => 
                           new_pc_value(20), inputs(12) => new_pc_value(19), 
                           inputs(13) => new_pc_value(18), inputs(14) => 
                           new_pc_value(17), inputs(15) => new_pc_value(16), 
                           inputs(16) => new_pc_value(15), inputs(17) => 
                           new_pc_value(14), inputs(18) => new_pc_value(13), 
                           inputs(19) => new_pc_value(12), inputs(20) => 
                           new_pc_value(11), inputs(21) => new_pc_value(10), 
                           inputs(22) => new_pc_value(9), inputs(23) => 
                           new_pc_value(8), inputs(24) => new_pc_value(7), 
                           inputs(25) => new_pc_value(6), inputs(26) => 
                           new_pc_value(5), inputs(27) => new_pc_value(4), 
                           inputs(28) => new_pc_value(3), inputs(29) => 
                           new_pc_value(2), inputs(30) => new_pc_value(1), 
                           inputs(31) => new_pc_value(0), inputs(32) => 
                           alu_output_val(31), inputs(33) => alu_output_val(30)
                           , inputs(34) => alu_output_val(29), inputs(35) => 
                           alu_output_val(28), inputs(36) => alu_output_val(27)
                           , inputs(37) => alu_output_val(26), inputs(38) => 
                           alu_output_val(25), inputs(39) => alu_output_val(24)
                           , inputs(40) => alu_output_val(23), inputs(41) => 
                           alu_output_val(22), inputs(42) => alu_output_val(21)
                           , inputs(43) => alu_output_val(20), inputs(44) => 
                           alu_output_val(19), inputs(45) => alu_output_val(18)
                           , inputs(46) => alu_output_val(17), inputs(47) => 
                           alu_output_val(16), inputs(48) => alu_output_val(15)
                           , inputs(49) => alu_output_val(14), inputs(50) => 
                           alu_output_val(13), inputs(51) => alu_output_val(12)
                           , inputs(52) => alu_output_val(11), inputs(53) => 
                           alu_output_val(10), inputs(54) => alu_output_val(9),
                           inputs(55) => alu_output_val(8), inputs(56) => 
                           alu_output_val(7), inputs(57) => alu_output_val(6), 
                           inputs(58) => alu_output_val(5), inputs(59) => 
                           alu_output_val(4), inputs(60) => alu_output_val(3), 
                           inputs(61) => alu_output_val(2), inputs(62) => 
                           alu_output_val(1), inputs(63) => alu_output_val(0), 
                           SEL => select_pc, Y(31) => new_pc_value_branch(31), 
                           Y(30) => new_pc_value_branch(30), Y(29) => 
                           new_pc_value_branch(29), Y(28) => 
                           new_pc_value_branch(28), Y(27) => 
                           new_pc_value_branch(27), Y(26) => 
                           new_pc_value_branch(26), Y(25) => 
                           new_pc_value_branch(25), Y(24) => 
                           new_pc_value_branch(24), Y(23) => 
                           new_pc_value_branch(23), Y(22) => 
                           new_pc_value_branch(22), Y(21) => 
                           new_pc_value_branch(21), Y(20) => 
                           new_pc_value_branch(20), Y(19) => 
                           new_pc_value_branch(19), Y(18) => 
                           new_pc_value_branch(18), Y(17) => 
                           new_pc_value_branch(17), Y(16) => 
                           new_pc_value_branch(16), Y(15) => 
                           new_pc_value_branch(15), Y(14) => 
                           new_pc_value_branch(14), Y(13) => 
                           new_pc_value_branch(13), Y(12) => 
                           new_pc_value_branch(12), Y(11) => 
                           new_pc_value_branch(11), Y(10) => 
                           new_pc_value_branch(10), Y(9) => 
                           new_pc_value_branch(9), Y(8) => 
                           new_pc_value_branch(8), Y(7) => 
                           new_pc_value_branch(7), Y(6) => 
                           new_pc_value_branch(6), Y(5) => 
                           new_pc_value_branch(5), Y(4) => 
                           new_pc_value_branch(4), Y(3) => 
                           new_pc_value_branch(3), Y(2) => 
                           new_pc_value_branch(2), Y(1) => 
                           new_pc_value_branch(1), Y(0) => 
                           new_pc_value_branch(0));
   lmd : reg_nbit_n32_8 port map( clk => clk, reset => n3, d(31) => 
                           data_ir_31_port, d(30) => data_ir_30_port, d(29) => 
                           data_ir_29_port, d(28) => data_ir_28_port, d(27) => 
                           data_ir_27_port, d(26) => data_ir_26_port, d(25) => 
                           data_ir_25_port, d(24) => data_ir_24_port, d(23) => 
                           data_ir_23_port, d(22) => data_ir_22_port, d(21) => 
                           data_ir_21_port, d(20) => data_ir_20_port, d(19) => 
                           data_ir_19_port, d(18) => data_ir_18_port, d(17) => 
                           data_ir_17_port, d(16) => data_ir_16_port, d(15) => 
                           data_ir_15_port, d(14) => data_ir_14_port, d(13) => 
                           data_ir_13_port, d(12) => data_ir_12_port, d(11) => 
                           data_ir_11_port, d(10) => data_ir_10_port, d(9) => 
                           data_ir_9_port, d(8) => data_ir_8_port, d(7) => 
                           data_ir_7_port, d(6) => data_ir_6_port, d(5) => 
                           data_ir_5_port, d(4) => data_ir_4_port, d(3) => 
                           data_ir_3_port, d(2) => data_ir_2_port, d(1) => 
                           data_ir_1_port, d(0) => data_ir_0_port, Q(31) => 
                           data_from_memory(31), Q(30) => data_from_memory(30),
                           Q(29) => data_from_memory(29), Q(28) => 
                           data_from_memory(28), Q(27) => data_from_memory(27),
                           Q(26) => data_from_memory(26), Q(25) => 
                           data_from_memory(25), Q(24) => data_from_memory(24),
                           Q(23) => data_from_memory(23), Q(22) => 
                           data_from_memory(22), Q(21) => data_from_memory(21),
                           Q(20) => data_from_memory(20), Q(19) => 
                           data_from_memory(19), Q(18) => data_from_memory(18),
                           Q(17) => data_from_memory(17), Q(16) => 
                           data_from_memory(16), Q(15) => data_from_memory(15),
                           Q(14) => data_from_memory(14), Q(13) => 
                           data_from_memory(13), Q(12) => data_from_memory(12),
                           Q(11) => data_from_memory(11), Q(10) => 
                           data_from_memory(10), Q(9) => data_from_memory(9), 
                           Q(8) => data_from_memory(8), Q(7) => 
                           data_from_memory(7), Q(6) => data_from_memory(6), 
                           Q(5) => data_from_memory(5), Q(4) => 
                           data_from_memory(4), Q(3) => data_from_memory(3), 
                           Q(2) => data_from_memory(2), Q(1) => 
                           data_from_memory(1), Q(0) => data_from_memory(0));
   delay_regg : reg_nbit_n32_7 port map( clk => clk, reset => n3, d(31) => 
                           alu_output_val(31), d(30) => alu_output_val(30), 
                           d(29) => alu_output_val(29), d(28) => 
                           alu_output_val(28), d(27) => alu_output_val(27), 
                           d(26) => alu_output_val(26), d(25) => 
                           alu_output_val(25), d(24) => alu_output_val(24), 
                           d(23) => alu_output_val(23), d(22) => 
                           alu_output_val(22), d(21) => alu_output_val(21), 
                           d(20) => alu_output_val(20), d(19) => 
                           alu_output_val(19), d(18) => alu_output_val(18), 
                           d(17) => alu_output_val(17), d(16) => 
                           alu_output_val(16), d(15) => alu_output_val(15), 
                           d(14) => alu_output_val(14), d(13) => 
                           alu_output_val(13), d(12) => alu_output_val(12), 
                           d(11) => alu_output_val(11), d(10) => 
                           alu_output_val(10), d(9) => alu_output_val(9), d(8) 
                           => alu_output_val(8), d(7) => alu_output_val(7), 
                           d(6) => alu_output_val(6), d(5) => alu_output_val(5)
                           , d(4) => alu_output_val(4), d(3) => 
                           alu_output_val(3), d(2) => alu_output_val(2), d(1) 
                           => alu_output_val(1), d(0) => alu_output_val(0), 
                           Q(31) => data_from_alu(31), Q(30) => 
                           data_from_alu(30), Q(29) => data_from_alu(29), Q(28)
                           => data_from_alu(28), Q(27) => data_from_alu(27), 
                           Q(26) => data_from_alu(26), Q(25) => 
                           data_from_alu(25), Q(24) => data_from_alu(24), Q(23)
                           => data_from_alu(23), Q(22) => data_from_alu(22), 
                           Q(21) => data_from_alu(21), Q(20) => 
                           data_from_alu(20), Q(19) => data_from_alu(19), Q(18)
                           => data_from_alu(18), Q(17) => data_from_alu(17), 
                           Q(16) => data_from_alu(16), Q(15) => 
                           data_from_alu(15), Q(14) => data_from_alu(14), Q(13)
                           => data_from_alu(13), Q(12) => data_from_alu(12), 
                           Q(11) => data_from_alu(11), Q(10) => 
                           data_from_alu(10), Q(9) => data_from_alu(9), Q(8) =>
                           data_from_alu(8), Q(7) => data_from_alu(7), Q(6) => 
                           data_from_alu(6), Q(5) => data_from_alu(5), Q(4) => 
                           data_from_alu(4), Q(3) => data_from_alu(3), Q(2) => 
                           data_from_alu(2), Q(1) => data_from_alu(1), Q(0) => 
                           data_from_alu(0));
   DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => value_to_mem(0), EN => n2, Z 
                           => DRAM_DATA(0));
   DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => value_to_mem(1), EN => n2, Z 
                           => DRAM_DATA(1));
   DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => value_to_mem(2), EN => n2, Z 
                           => DRAM_DATA(2));
   DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => value_to_mem(3), EN => n2, Z 
                           => DRAM_DATA(3));
   DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => value_to_mem(4), EN => n2, Z 
                           => DRAM_DATA(4));
   DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => value_to_mem(5), EN => n2, Z 
                           => DRAM_DATA(5));
   DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => value_to_mem(6), EN => n2, Z 
                           => DRAM_DATA(6));
   DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => value_to_mem(7), EN => n2, Z 
                           => DRAM_DATA(7));
   DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => value_to_mem(8), EN => n2, Z 
                           => DRAM_DATA(8));
   DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => value_to_mem(10), EN => n2, Z
                           => DRAM_DATA(10));
   DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => value_to_mem(11), EN => n2, Z
                           => DRAM_DATA(11));
   DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => value_to_mem(12), EN => n2, Z
                           => DRAM_DATA(12));
   DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => value_to_mem(13), EN => n2, Z
                           => DRAM_DATA(13));
   DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => value_to_mem(14), EN => n2, Z
                           => DRAM_DATA(14));
   DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => value_to_mem(15), EN => n2, Z
                           => DRAM_DATA(15));
   DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => value_to_mem(16), EN => n2, Z
                           => DRAM_DATA(16));
   DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => value_to_mem(17), EN => n2, Z
                           => DRAM_DATA(17));
   DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => value_to_mem(18), EN => n2, Z
                           => DRAM_DATA(18));
   DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => value_to_mem(19), EN => n2, Z
                           => DRAM_DATA(19));
   DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => value_to_mem(20), EN => n2, Z
                           => DRAM_DATA(20));
   DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => value_to_mem(21), EN => n2, Z
                           => DRAM_DATA(21));
   DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => value_to_mem(22), EN => n2, Z
                           => DRAM_DATA(22));
   DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => value_to_mem(23), EN => n2, Z
                           => DRAM_DATA(23));
   DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => value_to_mem(24), EN => n2, Z
                           => DRAM_DATA(24));
   DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => value_to_mem(25), EN => n2, Z
                           => DRAM_DATA(25));
   DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => value_to_mem(26), EN => n2, Z
                           => DRAM_DATA(26));
   DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => value_to_mem(27), EN => n2, Z
                           => DRAM_DATA(27));
   DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => value_to_mem(28), EN => n2, Z
                           => DRAM_DATA(28));
   DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => value_to_mem(29), EN => n2, Z
                           => DRAM_DATA(29));
   DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => value_to_mem(30), EN => n2, Z
                           => DRAM_DATA(30));
   DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => value_to_mem(31), EN => n2, Z
                           => DRAM_DATA(31));
   DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => value_to_mem(9), EN => n2, Z 
                           => DRAM_DATA(9));
   DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => alu_output_val(2), EN => n1
                           , Z => DRAM_ADDRESS_2_port);
   DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => alu_output_val(3), EN => n1
                           , Z => DRAM_ADDRESS_3_port);
   DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => alu_output_val(4), EN => n1
                           , Z => DRAM_ADDRESS_4_port);
   DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => alu_output_val(5), EN => n1
                           , Z => DRAM_ADDRESS_5_port);
   DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => alu_output_val(6), EN => n1
                           , Z => DRAM_ADDRESS_6_port);
   DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => alu_output_val(7), EN => n1
                           , Z => DRAM_ADDRESS_7_port);
   DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => alu_output_val(8), EN => n1
                           , Z => DRAM_ADDRESS_8_port);
   DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => alu_output_val(9), EN => n1
                           , Z => DRAM_ADDRESS_9_port);
   DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A => alu_output_val(10), EN => 
                           n1, Z => DRAM_ADDRESS_10_port);
   DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A => alu_output_val(11), EN => 
                           n1, Z => DRAM_ADDRESS_11_port);
   DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A => alu_output_val(12), EN => 
                           n1, Z => DRAM_ADDRESS_12_port);
   DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A => alu_output_val(13), EN => 
                           n1, Z => DRAM_ADDRESS_13_port);
   DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A => alu_output_val(14), EN => 
                           n1, Z => DRAM_ADDRESS_14_port);
   DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A => alu_output_val(15), EN => 
                           n1, Z => DRAM_ADDRESS_15_port);
   DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A => alu_output_val(16), EN => 
                           n1, Z => DRAM_ADDRESS_16_port);
   DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A => alu_output_val(17), EN => 
                           n1, Z => DRAM_ADDRESS_17_port);
   DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A => alu_output_val(18), EN => 
                           n1, Z => DRAM_ADDRESS_18_port);
   DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A => alu_output_val(19), EN => 
                           n1, Z => DRAM_ADDRESS_19_port);
   DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A => alu_output_val(20), EN => 
                           n1, Z => DRAM_ADDRESS_20_port);
   DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A => alu_output_val(21), EN => 
                           n1, Z => DRAM_ADDRESS_21_port);
   DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A => alu_output_val(22), EN => 
                           n1, Z => DRAM_ADDRESS_22_port);
   DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A => alu_output_val(23), EN => 
                           n1, Z => DRAM_ADDRESS_23_port);
   DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A => alu_output_val(24), EN => 
                           n1, Z => DRAM_ADDRESS_24_port);
   DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A => alu_output_val(25), EN => 
                           n1, Z => DRAM_ADDRESS_25_port);
   DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A => alu_output_val(26), EN => 
                           n1, Z => DRAM_ADDRESS_26_port);
   DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A => alu_output_val(27), EN => 
                           n1, Z => DRAM_ADDRESS_27_port);
   DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A => alu_output_val(28), EN => 
                           n1, Z => DRAM_ADDRESS_28_port);
   DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A => alu_output_val(29), EN => 
                           n1, Z => DRAM_ADDRESS_29_port);
   DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A => alu_output_val(30), EN => 
                           n1, Z => DRAM_ADDRESS_30_port);
   DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A => alu_output_val(31), EN => 
                           n1, Z => DRAM_ADDRESS_31_port);
   U2 : INV_X4 port map( A => rst, ZN => n3);
   U3 : INV_X2 port map( A => dram_enable_cu, ZN => n1);
   U4 : OR2_X2 port map( A1 => dram_r_nw_cu, A2 => n1, ZN => n2);
   U5 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           data_ir_9_port);
   U6 : AND2_X1 port map( A1 => DRAM_DATA(8), A2 => DRAM_READY, ZN => 
                           data_ir_8_port);
   U7 : AND2_X1 port map( A1 => DRAM_DATA(7), A2 => DRAM_READY, ZN => 
                           data_ir_7_port);
   U8 : AND2_X1 port map( A1 => DRAM_DATA(6), A2 => DRAM_READY, ZN => 
                           data_ir_6_port);
   U9 : AND2_X1 port map( A1 => DRAM_DATA(5), A2 => DRAM_READY, ZN => 
                           data_ir_5_port);
   U10 : AND2_X1 port map( A1 => DRAM_DATA(4), A2 => DRAM_READY, ZN => 
                           data_ir_4_port);
   U11 : AND2_X1 port map( A1 => DRAM_DATA(3), A2 => DRAM_READY, ZN => 
                           data_ir_3_port);
   U12 : AND2_X1 port map( A1 => DRAM_DATA(31), A2 => DRAM_READY, ZN => 
                           data_ir_31_port);
   U13 : AND2_X1 port map( A1 => DRAM_DATA(30), A2 => DRAM_READY, ZN => 
                           data_ir_30_port);
   U14 : AND2_X1 port map( A1 => DRAM_DATA(2), A2 => DRAM_READY, ZN => 
                           data_ir_2_port);
   U15 : AND2_X1 port map( A1 => DRAM_DATA(29), A2 => DRAM_READY, ZN => 
                           data_ir_29_port);
   U16 : AND2_X1 port map( A1 => DRAM_DATA(28), A2 => DRAM_READY, ZN => 
                           data_ir_28_port);
   U17 : AND2_X1 port map( A1 => DRAM_DATA(27), A2 => DRAM_READY, ZN => 
                           data_ir_27_port);
   U18 : AND2_X1 port map( A1 => DRAM_DATA(26), A2 => DRAM_READY, ZN => 
                           data_ir_26_port);
   U19 : AND2_X1 port map( A1 => DRAM_DATA(25), A2 => DRAM_READY, ZN => 
                           data_ir_25_port);
   U20 : AND2_X1 port map( A1 => DRAM_DATA(24), A2 => DRAM_READY, ZN => 
                           data_ir_24_port);
   U21 : AND2_X1 port map( A1 => DRAM_DATA(23), A2 => DRAM_READY, ZN => 
                           data_ir_23_port);
   U22 : AND2_X1 port map( A1 => DRAM_DATA(22), A2 => DRAM_READY, ZN => 
                           data_ir_22_port);
   U23 : AND2_X1 port map( A1 => DRAM_DATA(21), A2 => DRAM_READY, ZN => 
                           data_ir_21_port);
   U24 : AND2_X1 port map( A1 => DRAM_DATA(20), A2 => DRAM_READY, ZN => 
                           data_ir_20_port);
   U25 : AND2_X1 port map( A1 => DRAM_DATA(1), A2 => DRAM_READY, ZN => 
                           data_ir_1_port);
   U26 : AND2_X1 port map( A1 => DRAM_DATA(19), A2 => DRAM_READY, ZN => 
                           data_ir_19_port);
   U27 : AND2_X1 port map( A1 => DRAM_DATA(18), A2 => DRAM_READY, ZN => 
                           data_ir_18_port);
   U28 : AND2_X1 port map( A1 => DRAM_DATA(17), A2 => DRAM_READY, ZN => 
                           data_ir_17_port);
   U29 : AND2_X1 port map( A1 => DRAM_DATA(16), A2 => DRAM_READY, ZN => 
                           data_ir_16_port);
   U30 : AND2_X1 port map( A1 => DRAM_DATA(15), A2 => DRAM_READY, ZN => 
                           data_ir_15_port);
   U31 : AND2_X1 port map( A1 => DRAM_DATA(14), A2 => DRAM_READY, ZN => 
                           data_ir_14_port);
   U32 : AND2_X1 port map( A1 => DRAM_DATA(13), A2 => DRAM_READY, ZN => 
                           data_ir_13_port);
   U33 : AND2_X1 port map( A1 => DRAM_DATA(12), A2 => DRAM_READY, ZN => 
                           data_ir_12_port);
   U34 : AND2_X1 port map( A1 => DRAM_DATA(11), A2 => DRAM_READY, ZN => 
                           data_ir_11_port);
   U35 : AND2_X1 port map( A1 => DRAM_DATA(10), A2 => DRAM_READY, ZN => 
                           data_ir_10_port);
   U36 : AND2_X1 port map( A1 => DRAM_DATA(0), A2 => DRAM_READY, ZN => 
                           data_ir_0_port);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity execute_stage_N32_PC_SIZE32 is

   port( clk, rst : in std_logic;  val_a, val_b, val_immediate, 
         new_prog_counter_val_exe : in std_logic_vector (31 downto 0);  
         branch_condition : out std_logic;  prog_counter_forwaded, 
         alu_output_val, value_to_mem : out std_logic_vector (31 downto 0);  
         signed_notsigned : in std_logic;  alu_op_type : in std_logic_vector (3
         downto 0);  sel_val_a, sel_val_b, cin : in std_logic;  overflow, 
         zero_mul_detect, mul_exeception : out std_logic;  evaluate_branch : in
         std_logic_vector (1 downto 0));

end execute_stage_N32_PC_SIZE32;

architecture SYN_structural of execute_stage_N32_PC_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component reg_nbit_n32_9
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_10
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component general_alu_N32
      port( clk, rst : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX_zbit_nbit_N32_Z1_3
      port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX_zbit_nbit_N32_Z1_4
      port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n1
      port( clk, reset, d : in std_logic;  Q : out std_logic);
   end component;
   
   component check_branch_logic_N32
      port( input_val : in std_logic_vector (31 downto 0);  enable : in 
            std_logic;  decision : out std_logic);
   end component;
   
   signal evaluate_branch_enable, branch_taken_0_port, 
      branch_taken_reg_q_0_port, opa_31_port, opa_30_port, opa_29_port, 
      opa_28_port, opa_27_port, opa_26_port, opa_25_port, opa_24_port, 
      opa_23_port, opa_22_port, opa_21_port, opa_20_port, opa_19_port, 
      opa_18_port, opa_17_port, opa_16_port, opa_15_port, opa_14_port, 
      opa_13_port, opa_12_port, opa_11_port, opa_10_port, opa_9_port, 
      opa_8_port, opa_7_port, opa_6_port, opa_5_port, opa_4_port, opa_3_port, 
      opa_2_port, opa_1_port, opa_0_port, opb_31_port, opb_30_port, opb_29_port
      , opb_28_port, opb_27_port, opb_26_port, opb_25_port, opb_24_port, 
      opb_23_port, opb_22_port, opb_21_port, opb_20_port, opb_19_port, 
      opb_18_port, opb_17_port, opb_16_port, opb_15_port, opb_14_port, 
      opb_13_port, opb_12_port, opb_11_port, opb_10_port, opb_9_port, 
      opb_8_port, opb_7_port, opb_6_port, opb_5_port, opb_4_port, opb_3_port, 
      opb_2_port, opb_1_port, opb_0_port, alu_op_type_i_3_port, 
      alu_op_type_i_1_port, alu_op_type_i_0_port, alu_out_31_port, 
      alu_out_30_port, alu_out_29_port, alu_out_28_port, alu_out_27_port, 
      alu_out_26_port, alu_out_25_port, alu_out_24_port, alu_out_23_port, 
      alu_out_22_port, alu_out_21_port, alu_out_20_port, alu_out_19_port, 
      alu_out_18_port, alu_out_17_port, alu_out_16_port, alu_out_15_port, 
      alu_out_14_port, alu_out_13_port, alu_out_12_port, alu_out_11_port, 
      alu_out_10_port, alu_out_9_port, alu_out_8_port, alu_out_7_port, 
      alu_out_6_port, alu_out_5_port, alu_out_4_port, alu_out_3_port, 
      alu_out_2_port, alu_out_1_port, alu_out_0_port, n1, n2, n3, n4, n5, n6, 
      n7, n8 : std_logic;

begin
   prog_counter_forwaded <= ( new_prog_counter_val_exe(31), 
      new_prog_counter_val_exe(30), new_prog_counter_val_exe(29), 
      new_prog_counter_val_exe(28), new_prog_counter_val_exe(27), 
      new_prog_counter_val_exe(26), new_prog_counter_val_exe(25), 
      new_prog_counter_val_exe(24), new_prog_counter_val_exe(23), 
      new_prog_counter_val_exe(22), new_prog_counter_val_exe(21), 
      new_prog_counter_val_exe(20), new_prog_counter_val_exe(19), 
      new_prog_counter_val_exe(18), new_prog_counter_val_exe(17), 
      new_prog_counter_val_exe(16), new_prog_counter_val_exe(15), 
      new_prog_counter_val_exe(14), new_prog_counter_val_exe(13), 
      new_prog_counter_val_exe(12), new_prog_counter_val_exe(11), 
      new_prog_counter_val_exe(10), new_prog_counter_val_exe(9), 
      new_prog_counter_val_exe(8), new_prog_counter_val_exe(7), 
      new_prog_counter_val_exe(6), new_prog_counter_val_exe(5), 
      new_prog_counter_val_exe(4), new_prog_counter_val_exe(3), 
      new_prog_counter_val_exe(2), new_prog_counter_val_exe(1), 
      new_prog_counter_val_exe(0) );
   
   check_branch_logic_i : check_branch_logic_N32 port map( input_val(31) => 
                           val_a(31), input_val(30) => val_a(30), input_val(29)
                           => val_a(29), input_val(28) => val_a(28), 
                           input_val(27) => val_a(27), input_val(26) => 
                           val_a(26), input_val(25) => val_a(25), input_val(24)
                           => val_a(24), input_val(23) => val_a(23), 
                           input_val(22) => val_a(22), input_val(21) => 
                           val_a(21), input_val(20) => val_a(20), input_val(19)
                           => val_a(19), input_val(18) => val_a(18), 
                           input_val(17) => val_a(17), input_val(16) => 
                           val_a(16), input_val(15) => val_a(15), input_val(14)
                           => val_a(14), input_val(13) => val_a(13), 
                           input_val(12) => val_a(12), input_val(11) => 
                           val_a(11), input_val(10) => val_a(10), input_val(9) 
                           => val_a(9), input_val(8) => val_a(8), input_val(7) 
                           => val_a(7), input_val(6) => val_a(6), input_val(5) 
                           => val_a(5), input_val(4) => val_a(4), input_val(3) 
                           => val_a(3), input_val(2) => val_a(2), input_val(1) 
                           => val_a(1), input_val(0) => val_a(0), enable => 
                           evaluate_branch_enable, decision => 
                           branch_taken_0_port);
   condition_delay_reg : reg_nbit_n1 port map( clk => clk, reset => n8, d => 
                           branch_taken_reg_q_0_port, Q => branch_condition);
   alu_opa : MUX_zbit_nbit_N32_Z1_4 port map( inputs(0) => val_a(31), inputs(1)
                           => val_a(30), inputs(2) => val_a(29), inputs(3) => 
                           val_a(28), inputs(4) => val_a(27), inputs(5) => 
                           val_a(26), inputs(6) => val_a(25), inputs(7) => 
                           val_a(24), inputs(8) => val_a(23), inputs(9) => 
                           val_a(22), inputs(10) => val_a(21), inputs(11) => 
                           val_a(20), inputs(12) => val_a(19), inputs(13) => 
                           val_a(18), inputs(14) => val_a(17), inputs(15) => 
                           val_a(16), inputs(16) => val_a(15), inputs(17) => 
                           val_a(14), inputs(18) => val_a(13), inputs(19) => 
                           val_a(12), inputs(20) => val_a(11), inputs(21) => 
                           val_a(10), inputs(22) => val_a(9), inputs(23) => 
                           val_a(8), inputs(24) => val_a(7), inputs(25) => 
                           val_a(6), inputs(26) => val_a(5), inputs(27) => 
                           val_a(4), inputs(28) => val_a(3), inputs(29) => 
                           val_a(2), inputs(30) => val_a(1), inputs(31) => 
                           val_a(0), inputs(32) => new_prog_counter_val_exe(31)
                           , inputs(33) => new_prog_counter_val_exe(30), 
                           inputs(34) => new_prog_counter_val_exe(29), 
                           inputs(35) => new_prog_counter_val_exe(28), 
                           inputs(36) => new_prog_counter_val_exe(27), 
                           inputs(37) => new_prog_counter_val_exe(26), 
                           inputs(38) => new_prog_counter_val_exe(25), 
                           inputs(39) => new_prog_counter_val_exe(24), 
                           inputs(40) => new_prog_counter_val_exe(23), 
                           inputs(41) => new_prog_counter_val_exe(22), 
                           inputs(42) => new_prog_counter_val_exe(21), 
                           inputs(43) => new_prog_counter_val_exe(20), 
                           inputs(44) => new_prog_counter_val_exe(19), 
                           inputs(45) => new_prog_counter_val_exe(18), 
                           inputs(46) => new_prog_counter_val_exe(17), 
                           inputs(47) => new_prog_counter_val_exe(16), 
                           inputs(48) => new_prog_counter_val_exe(15), 
                           inputs(49) => new_prog_counter_val_exe(14), 
                           inputs(50) => new_prog_counter_val_exe(13), 
                           inputs(51) => new_prog_counter_val_exe(12), 
                           inputs(52) => new_prog_counter_val_exe(11), 
                           inputs(53) => new_prog_counter_val_exe(10), 
                           inputs(54) => new_prog_counter_val_exe(9), 
                           inputs(55) => new_prog_counter_val_exe(8), 
                           inputs(56) => new_prog_counter_val_exe(7), 
                           inputs(57) => new_prog_counter_val_exe(6), 
                           inputs(58) => new_prog_counter_val_exe(5), 
                           inputs(59) => new_prog_counter_val_exe(4), 
                           inputs(60) => new_prog_counter_val_exe(3), 
                           inputs(61) => new_prog_counter_val_exe(2), 
                           inputs(62) => new_prog_counter_val_exe(1), 
                           inputs(63) => new_prog_counter_val_exe(0), SEL => 
                           sel_val_a, Y(31) => opa_31_port, Y(30) => 
                           opa_30_port, Y(29) => opa_29_port, Y(28) => 
                           opa_28_port, Y(27) => opa_27_port, Y(26) => 
                           opa_26_port, Y(25) => opa_25_port, Y(24) => 
                           opa_24_port, Y(23) => opa_23_port, Y(22) => 
                           opa_22_port, Y(21) => opa_21_port, Y(20) => 
                           opa_20_port, Y(19) => opa_19_port, Y(18) => 
                           opa_18_port, Y(17) => opa_17_port, Y(16) => 
                           opa_16_port, Y(15) => opa_15_port, Y(14) => 
                           opa_14_port, Y(13) => opa_13_port, Y(12) => 
                           opa_12_port, Y(11) => opa_11_port, Y(10) => 
                           opa_10_port, Y(9) => opa_9_port, Y(8) => opa_8_port,
                           Y(7) => opa_7_port, Y(6) => opa_6_port, Y(5) => 
                           opa_5_port, Y(4) => opa_4_port, Y(3) => opa_3_port, 
                           Y(2) => opa_2_port, Y(1) => opa_1_port, Y(0) => 
                           opa_0_port);
   alu_opb : MUX_zbit_nbit_N32_Z1_3 port map( inputs(0) => val_b(31), inputs(1)
                           => val_b(30), inputs(2) => val_b(29), inputs(3) => 
                           val_b(28), inputs(4) => val_b(27), inputs(5) => 
                           val_b(26), inputs(6) => val_b(25), inputs(7) => 
                           val_b(24), inputs(8) => val_b(23), inputs(9) => 
                           val_b(22), inputs(10) => val_b(21), inputs(11) => 
                           val_b(20), inputs(12) => val_b(19), inputs(13) => 
                           val_b(18), inputs(14) => val_b(17), inputs(15) => 
                           val_b(16), inputs(16) => val_b(15), inputs(17) => 
                           val_b(14), inputs(18) => val_b(13), inputs(19) => 
                           val_b(12), inputs(20) => val_b(11), inputs(21) => 
                           val_b(10), inputs(22) => val_b(9), inputs(23) => 
                           val_b(8), inputs(24) => val_b(7), inputs(25) => 
                           val_b(6), inputs(26) => val_b(5), inputs(27) => 
                           val_b(4), inputs(28) => val_b(3), inputs(29) => 
                           val_b(2), inputs(30) => val_b(1), inputs(31) => 
                           val_b(0), inputs(32) => val_immediate(31), 
                           inputs(33) => val_immediate(30), inputs(34) => 
                           val_immediate(29), inputs(35) => val_immediate(28), 
                           inputs(36) => val_immediate(27), inputs(37) => 
                           val_immediate(26), inputs(38) => val_immediate(25), 
                           inputs(39) => val_immediate(24), inputs(40) => 
                           val_immediate(23), inputs(41) => val_immediate(22), 
                           inputs(42) => val_immediate(21), inputs(43) => 
                           val_immediate(20), inputs(44) => val_immediate(19), 
                           inputs(45) => val_immediate(18), inputs(46) => 
                           val_immediate(17), inputs(47) => val_immediate(16), 
                           inputs(48) => val_immediate(15), inputs(49) => 
                           val_immediate(14), inputs(50) => val_immediate(13), 
                           inputs(51) => val_immediate(12), inputs(52) => 
                           val_immediate(11), inputs(53) => val_immediate(10), 
                           inputs(54) => val_immediate(9), inputs(55) => 
                           val_immediate(8), inputs(56) => val_immediate(7), 
                           inputs(57) => val_immediate(6), inputs(58) => 
                           val_immediate(5), inputs(59) => val_immediate(4), 
                           inputs(60) => val_immediate(3), inputs(61) => 
                           val_immediate(2), inputs(62) => val_immediate(1), 
                           inputs(63) => val_immediate(0), SEL => sel_val_b, 
                           Y(31) => opb_31_port, Y(30) => opb_30_port, Y(29) =>
                           opb_29_port, Y(28) => opb_28_port, Y(27) => 
                           opb_27_port, Y(26) => opb_26_port, Y(25) => 
                           opb_25_port, Y(24) => opb_24_port, Y(23) => 
                           opb_23_port, Y(22) => opb_22_port, Y(21) => 
                           opb_21_port, Y(20) => opb_20_port, Y(19) => 
                           opb_19_port, Y(18) => opb_18_port, Y(17) => 
                           opb_17_port, Y(16) => opb_16_port, Y(15) => 
                           opb_15_port, Y(14) => opb_14_port, Y(13) => 
                           opb_13_port, Y(12) => opb_12_port, Y(11) => 
                           opb_11_port, Y(10) => opb_10_port, Y(9) => 
                           opb_9_port, Y(8) => opb_8_port, Y(7) => opb_7_port, 
                           Y(6) => opb_6_port, Y(5) => opb_5_port, Y(4) => 
                           opb_4_port, Y(3) => opb_3_port, Y(2) => opb_2_port, 
                           Y(1) => opb_1_port, Y(0) => opb_0_port);
   general_alu_i : general_alu_N32 port map( clk => clk, rst => n8, 
                           zero_mul_detect => zero_mul_detect, mul_exeception 
                           => mul_exeception, FUNC(0) => alu_op_type_i_3_port, 
                           FUNC(1) => n7, FUNC(2) => alu_op_type_i_1_port, 
                           FUNC(3) => alu_op_type_i_0_port, DATA1(31) => 
                           opa_31_port, DATA1(30) => opa_30_port, DATA1(29) => 
                           opa_29_port, DATA1(28) => opa_28_port, DATA1(27) => 
                           opa_27_port, DATA1(26) => opa_26_port, DATA1(25) => 
                           opa_25_port, DATA1(24) => opa_24_port, DATA1(23) => 
                           opa_23_port, DATA1(22) => opa_22_port, DATA1(21) => 
                           opa_21_port, DATA1(20) => opa_20_port, DATA1(19) => 
                           opa_19_port, DATA1(18) => opa_18_port, DATA1(17) => 
                           opa_17_port, DATA1(16) => opa_16_port, DATA1(15) => 
                           opa_15_port, DATA1(14) => opa_14_port, DATA1(13) => 
                           opa_13_port, DATA1(12) => opa_12_port, DATA1(11) => 
                           opa_11_port, DATA1(10) => opa_10_port, DATA1(9) => 
                           opa_9_port, DATA1(8) => opa_8_port, DATA1(7) => 
                           opa_7_port, DATA1(6) => opa_6_port, DATA1(5) => 
                           opa_5_port, DATA1(4) => opa_4_port, DATA1(3) => 
                           opa_3_port, DATA1(2) => opa_2_port, DATA1(1) => 
                           opa_1_port, DATA1(0) => opa_0_port, DATA2(31) => 
                           opb_31_port, DATA2(30) => opb_30_port, DATA2(29) => 
                           opb_29_port, DATA2(28) => opb_28_port, DATA2(27) => 
                           opb_27_port, DATA2(26) => opb_26_port, DATA2(25) => 
                           opb_25_port, DATA2(24) => opb_24_port, DATA2(23) => 
                           opb_23_port, DATA2(22) => opb_22_port, DATA2(21) => 
                           opb_21_port, DATA2(20) => opb_20_port, DATA2(19) => 
                           opb_19_port, DATA2(18) => opb_18_port, DATA2(17) => 
                           opb_17_port, DATA2(16) => opb_16_port, DATA2(15) => 
                           opb_15_port, DATA2(14) => opb_14_port, DATA2(13) => 
                           opb_13_port, DATA2(12) => opb_12_port, DATA2(11) => 
                           opb_11_port, DATA2(10) => opb_10_port, DATA2(9) => 
                           opb_9_port, DATA2(8) => opb_8_port, DATA2(7) => 
                           opb_7_port, DATA2(6) => opb_6_port, DATA2(5) => 
                           opb_5_port, DATA2(4) => opb_4_port, DATA2(3) => 
                           opb_3_port, DATA2(2) => opb_2_port, DATA2(1) => 
                           opb_1_port, DATA2(0) => opb_0_port, cin => cin, 
                           signed_notsigned => signed_notsigned, overflow => 
                           overflow, OUTALU(31) => alu_out_31_port, OUTALU(30) 
                           => alu_out_30_port, OUTALU(29) => alu_out_29_port, 
                           OUTALU(28) => alu_out_28_port, OUTALU(27) => 
                           alu_out_27_port, OUTALU(26) => alu_out_26_port, 
                           OUTALU(25) => alu_out_25_port, OUTALU(24) => 
                           alu_out_24_port, OUTALU(23) => alu_out_23_port, 
                           OUTALU(22) => alu_out_22_port, OUTALU(21) => 
                           alu_out_21_port, OUTALU(20) => alu_out_20_port, 
                           OUTALU(19) => alu_out_19_port, OUTALU(18) => 
                           alu_out_18_port, OUTALU(17) => alu_out_17_port, 
                           OUTALU(16) => alu_out_16_port, OUTALU(15) => 
                           alu_out_15_port, OUTALU(14) => alu_out_14_port, 
                           OUTALU(13) => alu_out_13_port, OUTALU(12) => 
                           alu_out_12_port, OUTALU(11) => alu_out_11_port, 
                           OUTALU(10) => alu_out_10_port, OUTALU(9) => 
                           alu_out_9_port, OUTALU(8) => alu_out_8_port, 
                           OUTALU(7) => alu_out_7_port, OUTALU(6) => 
                           alu_out_6_port, OUTALU(5) => alu_out_5_port, 
                           OUTALU(4) => alu_out_4_port, OUTALU(3) => 
                           alu_out_3_port, OUTALU(2) => alu_out_2_port, 
                           OUTALU(1) => alu_out_1_port, OUTALU(0) => 
                           alu_out_0_port);
   alu_reg_out : reg_nbit_n32_10 port map( clk => clk, reset => n8, d(31) => 
                           alu_out_31_port, d(30) => alu_out_30_port, d(29) => 
                           alu_out_29_port, d(28) => alu_out_28_port, d(27) => 
                           alu_out_27_port, d(26) => alu_out_26_port, d(25) => 
                           alu_out_25_port, d(24) => alu_out_24_port, d(23) => 
                           alu_out_23_port, d(22) => alu_out_22_port, d(21) => 
                           alu_out_21_port, d(20) => alu_out_20_port, d(19) => 
                           alu_out_19_port, d(18) => alu_out_18_port, d(17) => 
                           alu_out_17_port, d(16) => alu_out_16_port, d(15) => 
                           alu_out_15_port, d(14) => alu_out_14_port, d(13) => 
                           alu_out_13_port, d(12) => alu_out_12_port, d(11) => 
                           alu_out_11_port, d(10) => alu_out_10_port, d(9) => 
                           alu_out_9_port, d(8) => alu_out_8_port, d(7) => 
                           alu_out_7_port, d(6) => alu_out_6_port, d(5) => 
                           alu_out_5_port, d(4) => alu_out_4_port, d(3) => 
                           alu_out_3_port, d(2) => alu_out_2_port, d(1) => 
                           alu_out_1_port, d(0) => alu_out_0_port, Q(31) => 
                           alu_output_val(31), Q(30) => alu_output_val(30), 
                           Q(29) => alu_output_val(29), Q(28) => 
                           alu_output_val(28), Q(27) => alu_output_val(27), 
                           Q(26) => alu_output_val(26), Q(25) => 
                           alu_output_val(25), Q(24) => alu_output_val(24), 
                           Q(23) => alu_output_val(23), Q(22) => 
                           alu_output_val(22), Q(21) => alu_output_val(21), 
                           Q(20) => alu_output_val(20), Q(19) => 
                           alu_output_val(19), Q(18) => alu_output_val(18), 
                           Q(17) => alu_output_val(17), Q(16) => 
                           alu_output_val(16), Q(15) => alu_output_val(15), 
                           Q(14) => alu_output_val(14), Q(13) => 
                           alu_output_val(13), Q(12) => alu_output_val(12), 
                           Q(11) => alu_output_val(11), Q(10) => 
                           alu_output_val(10), Q(9) => alu_output_val(9), Q(8) 
                           => alu_output_val(8), Q(7) => alu_output_val(7), 
                           Q(6) => alu_output_val(6), Q(5) => alu_output_val(5)
                           , Q(4) => alu_output_val(4), Q(3) => 
                           alu_output_val(3), Q(2) => alu_output_val(2), Q(1) 
                           => alu_output_val(1), Q(0) => alu_output_val(0));
   reg_del_b : reg_nbit_n32_9 port map( clk => clk, reset => n8, d(31) => 
                           val_b(31), d(30) => val_b(30), d(29) => val_b(29), 
                           d(28) => val_b(28), d(27) => val_b(27), d(26) => 
                           val_b(26), d(25) => val_b(25), d(24) => val_b(24), 
                           d(23) => val_b(23), d(22) => val_b(22), d(21) => 
                           val_b(21), d(20) => val_b(20), d(19) => val_b(19), 
                           d(18) => val_b(18), d(17) => val_b(17), d(16) => 
                           val_b(16), d(15) => val_b(15), d(14) => val_b(14), 
                           d(13) => val_b(13), d(12) => val_b(12), d(11) => 
                           val_b(11), d(10) => val_b(10), d(9) => val_b(9), 
                           d(8) => val_b(8), d(7) => val_b(7), d(6) => val_b(6)
                           , d(5) => val_b(5), d(4) => val_b(4), d(3) => 
                           val_b(3), d(2) => val_b(2), d(1) => val_b(1), d(0) 
                           => val_b(0), Q(31) => value_to_mem(31), Q(30) => 
                           value_to_mem(30), Q(29) => value_to_mem(29), Q(28) 
                           => value_to_mem(28), Q(27) => value_to_mem(27), 
                           Q(26) => value_to_mem(26), Q(25) => value_to_mem(25)
                           , Q(24) => value_to_mem(24), Q(23) => 
                           value_to_mem(23), Q(22) => value_to_mem(22), Q(21) 
                           => value_to_mem(21), Q(20) => value_to_mem(20), 
                           Q(19) => value_to_mem(19), Q(18) => value_to_mem(18)
                           , Q(17) => value_to_mem(17), Q(16) => 
                           value_to_mem(16), Q(15) => value_to_mem(15), Q(14) 
                           => value_to_mem(14), Q(13) => value_to_mem(13), 
                           Q(12) => value_to_mem(12), Q(11) => value_to_mem(11)
                           , Q(10) => value_to_mem(10), Q(9) => value_to_mem(9)
                           , Q(8) => value_to_mem(8), Q(7) => value_to_mem(7), 
                           Q(6) => value_to_mem(6), Q(5) => value_to_mem(5), 
                           Q(4) => value_to_mem(4), Q(3) => value_to_mem(3), 
                           Q(2) => value_to_mem(2), Q(1) => value_to_mem(1), 
                           Q(0) => value_to_mem(0));
   U3 : NOR2_X1 port map( A1 => alu_op_type(3), A2 => n1, ZN => n7);
   U4 : INV_X1 port map( A => rst, ZN => n8);
   U5 : OR2_X1 port map( A1 => evaluate_branch(0), A2 => evaluate_branch(1), ZN
                           => evaluate_branch_enable);
   U6 : XOR2_X1 port map( A => evaluate_branch(1), B => branch_taken_0_port, Z 
                           => branch_taken_reg_q_0_port);
   U7 : AOI211_X1 port map( C1 => alu_op_type(1), C2 => alu_op_type(0), A => n2
                           , B => alu_op_type(2), ZN => alu_op_type_i_3_port);
   U8 : NOR2_X1 port map( A1 => n3, A2 => n4, ZN => alu_op_type_i_1_port);
   U9 : AOI21_X1 port map( B1 => n5, B2 => n1, A => n2, ZN => n3);
   U10 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => alu_op_type_i_0_port);
   U11 : INV_X1 port map( A => alu_op_type(0), ZN => n5);
   U12 : AOI21_X1 port map( B1 => n4, B2 => n1, A => n2, ZN => n6);
   U13 : INV_X1 port map( A => alu_op_type(3), ZN => n2);
   U14 : INV_X1 port map( A => alu_op_type(2), ZN => n1);
   U15 : INV_X1 port map( A => alu_op_type(1), ZN => n4);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity decode_stage_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 is

   port( clk, rst : in std_logic;  new_prog_counter_val, instruction_reg : in 
         std_logic_vector (31 downto 0);  val_a, new_prog_counter_val_exe, 
         val_b, val_immediate : out std_logic_vector (31 downto 0);  
         update_reg_value : in std_logic_vector (31 downto 0);  enable_rf, 
         read_rf_p1, read_rf_p2, write_rf, rtype_itypen, jump_sext, 
         compute_sext : in std_logic);

end decode_stage_N32_RF_REGS32_IR_SIZE32_PC_SIZE32;

architecture SYN_structural of decode_stage_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component reg_nbit_n33_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (32 downto 0); 
            Q : out std_logic_vector (32 downto 0));
   end component;
   
   component reg_nbit_n33_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (32 downto 0); 
            Q : out std_logic_vector (32 downto 0));
   end component;
   
   component reg_nbit_n32_11
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX_zbit_nbit_N32_Z1_0
      port( inputs : in std_logic_vector (0 to 63);  SEL : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component sign_extension_N32_STARTING_BIT26
      port( val_to_exetend : in std_logic_vector (25 downto 0);  enable : in 
            std_logic;  extended_val : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_extension_N32_STARTING_BIT16
      port( val_to_exetend : in std_logic_vector (15 downto 0);  enable : in 
            std_logic;  extended_val : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_12
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_13
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component reg_nbit_n5_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_nbit_n5_2
      port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_nbit_n5_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (4 downto 0);  
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   signal enable_sign_extension_logic, del_reg_wb_1_4_port, del_reg_wb_1_3_port
      , del_reg_wb_1_2_port, del_reg_wb_1_1_port, del_reg_wb_1_0_port, 
      del_reg_wb_2_4_port, del_reg_wb_2_3_port, del_reg_wb_2_2_port, 
      del_reg_wb_2_1_port, del_reg_wb_2_0_port, address_rf_write_4_port, 
      address_rf_write_3_port, address_rf_write_2_port, address_rf_write_1_port
      , address_rf_write_0_port, enable_rf_i, val_reg_a_i_31_port, 
      val_reg_a_i_30_port, val_reg_a_i_29_port, val_reg_a_i_28_port, 
      val_reg_a_i_27_port, val_reg_a_i_26_port, val_reg_a_i_25_port, 
      val_reg_a_i_24_port, val_reg_a_i_23_port, val_reg_a_i_22_port, 
      val_reg_a_i_21_port, val_reg_a_i_20_port, val_reg_a_i_19_port, 
      val_reg_a_i_18_port, val_reg_a_i_17_port, val_reg_a_i_16_port, 
      val_reg_a_i_15_port, val_reg_a_i_14_port, val_reg_a_i_13_port, 
      val_reg_a_i_12_port, val_reg_a_i_11_port, val_reg_a_i_10_port, 
      val_reg_a_i_9_port, val_reg_a_i_8_port, val_reg_a_i_7_port, 
      val_reg_a_i_6_port, val_reg_a_i_5_port, val_reg_a_i_4_port, 
      val_reg_a_i_3_port, val_reg_a_i_2_port, val_reg_a_i_1_port, 
      val_reg_a_i_0_port, val_reg_b_i_31_port, val_reg_b_i_30_port, 
      val_reg_b_i_29_port, val_reg_b_i_28_port, val_reg_b_i_27_port, 
      val_reg_b_i_26_port, val_reg_b_i_25_port, val_reg_b_i_24_port, 
      val_reg_b_i_23_port, val_reg_b_i_22_port, val_reg_b_i_21_port, 
      val_reg_b_i_20_port, val_reg_b_i_19_port, val_reg_b_i_18_port, 
      val_reg_b_i_17_port, val_reg_b_i_16_port, val_reg_b_i_15_port, 
      val_reg_b_i_14_port, val_reg_b_i_13_port, val_reg_b_i_12_port, 
      val_reg_b_i_11_port, val_reg_b_i_10_port, val_reg_b_i_9_port, 
      val_reg_b_i_8_port, val_reg_b_i_7_port, val_reg_b_i_6_port, 
      val_reg_b_i_5_port, val_reg_b_i_4_port, val_reg_b_i_3_port, 
      val_reg_b_i_2_port, val_reg_b_i_1_port, val_reg_b_i_0_port, 
      val_reg_immediate_i_31_port, val_reg_immediate_i_30_port, 
      val_reg_immediate_i_29_port, val_reg_immediate_i_28_port, 
      val_reg_immediate_i_27_port, val_reg_immediate_i_26_port, 
      val_reg_immediate_i_25_port, val_reg_immediate_i_24_port, 
      val_reg_immediate_i_23_port, val_reg_immediate_i_22_port, 
      val_reg_immediate_i_21_port, val_reg_immediate_i_20_port, 
      val_reg_immediate_i_19_port, val_reg_immediate_i_18_port, 
      val_reg_immediate_i_17_port, val_reg_immediate_i_16_port, 
      val_reg_immediate_i_15_port, val_reg_immediate_i_14_port, 
      val_reg_immediate_i_13_port, val_reg_immediate_i_12_port, 
      val_reg_immediate_i_11_port, val_reg_immediate_i_10_port, 
      val_reg_immediate_i_9_port, val_reg_immediate_i_8_port, 
      val_reg_immediate_i_7_port, val_reg_immediate_i_6_port, 
      val_reg_immediate_i_5_port, val_reg_immediate_i_4_port, 
      val_reg_immediate_i_3_port, val_reg_immediate_i_2_port, 
      val_reg_immediate_i_1_port, val_reg_immediate_i_0_port, 
      val_reg_immediate_j_31_port, val_reg_immediate_j_30_port, 
      val_reg_immediate_j_29_port, val_reg_immediate_j_28_port, 
      val_reg_immediate_j_27_port, val_reg_immediate_j_26_port, 
      val_reg_immediate_j_25_port, val_reg_immediate_j_24_port, 
      val_reg_immediate_j_23_port, val_reg_immediate_j_22_port, 
      val_reg_immediate_j_21_port, val_reg_immediate_j_20_port, 
      val_reg_immediate_j_19_port, val_reg_immediate_j_18_port, 
      val_reg_immediate_j_17_port, val_reg_immediate_j_16_port, 
      val_reg_immediate_j_15_port, val_reg_immediate_j_14_port, 
      val_reg_immediate_j_13_port, val_reg_immediate_j_12_port, 
      val_reg_immediate_j_11_port, val_reg_immediate_j_10_port, 
      val_reg_immediate_j_9_port, val_reg_immediate_j_8_port, 
      val_reg_immediate_j_7_port, val_reg_immediate_j_6_port, 
      val_reg_immediate_j_5_port, val_reg_immediate_j_4_port, 
      val_reg_immediate_j_3_port, val_reg_immediate_j_2_port, 
      val_reg_immediate_j_1_port, val_reg_immediate_j_0_port, 
      val_reg_immediate_31_port, val_reg_immediate_30_port, 
      val_reg_immediate_29_port, val_reg_immediate_28_port, 
      val_reg_immediate_27_port, val_reg_immediate_26_port, 
      val_reg_immediate_25_port, val_reg_immediate_24_port, 
      val_reg_immediate_23_port, val_reg_immediate_22_port, 
      val_reg_immediate_21_port, val_reg_immediate_20_port, 
      val_reg_immediate_19_port, val_reg_immediate_18_port, 
      val_reg_immediate_17_port, val_reg_immediate_16_port, 
      val_reg_immediate_15_port, val_reg_immediate_14_port, 
      val_reg_immediate_13_port, val_reg_immediate_12_port, 
      val_reg_immediate_11_port, val_reg_immediate_10_port, 
      val_reg_immediate_9_port, val_reg_immediate_8_port, 
      val_reg_immediate_7_port, val_reg_immediate_6_port, 
      val_reg_immediate_5_port, val_reg_immediate_4_port, 
      val_reg_immediate_3_port, val_reg_immediate_2_port, 
      val_reg_immediate_1_port, val_reg_immediate_0_port, clk_immediate, 
      pc_delay2_32_port, pc_delay2_31_port, pc_delay2_30_port, 
      pc_delay2_29_port, pc_delay2_28_port, pc_delay2_27_port, 
      pc_delay2_26_port, pc_delay2_25_port, pc_delay2_24_port, 
      pc_delay2_23_port, pc_delay2_22_port, pc_delay2_21_port, 
      pc_delay2_20_port, pc_delay2_19_port, pc_delay2_18_port, 
      pc_delay2_17_port, pc_delay2_16_port, pc_delay2_15_port, 
      pc_delay2_14_port, pc_delay2_13_port, pc_delay2_12_port, 
      pc_delay2_11_port, pc_delay2_10_port, pc_delay2_9_port, pc_delay2_8_port,
      pc_delay2_7_port, pc_delay2_6_port, pc_delay2_5_port, pc_delay2_4_port, 
      pc_delay2_3_port, pc_delay2_2_port, pc_delay2_1_port, pc_delay2_0_port, 
      pc_delay3_32_port, pc_delay3_31_port, pc_delay3_30_port, 
      pc_delay3_29_port, pc_delay3_28_port, pc_delay3_27_port, 
      pc_delay3_26_port, pc_delay3_25_port, pc_delay3_24_port, 
      pc_delay3_23_port, pc_delay3_22_port, pc_delay3_21_port, 
      pc_delay3_20_port, pc_delay3_19_port, pc_delay3_18_port, 
      pc_delay3_17_port, pc_delay3_16_port, pc_delay3_15_port, 
      pc_delay3_14_port, pc_delay3_13_port, pc_delay3_12_port, 
      pc_delay3_11_port, pc_delay3_10_port, pc_delay3_9_port, pc_delay3_8_port,
      pc_delay3_7_port, pc_delay3_6_port, pc_delay3_5_port, pc_delay3_4_port, 
      pc_delay3_3_port, pc_delay3_2_port, pc_delay3_1_port, pc_delay3_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n76, n77, 
      n78, n79, n80, n81, n82 : std_logic;

begin
   
   delay_reg_wb_1 : reg_nbit_n5_0 port map( clk => n2, reset => n1, d(4) => n80
                           , d(3) => n79, d(2) => n78, d(1) => n77, d(0) => n76
                           , Q(4) => del_reg_wb_1_4_port, Q(3) => 
                           del_reg_wb_1_3_port, Q(2) => del_reg_wb_1_2_port, 
                           Q(1) => del_reg_wb_1_1_port, Q(0) => 
                           del_reg_wb_1_0_port);
   delay_reg_wb_2 : reg_nbit_n5_2 port map( clk => n2, reset => n1, d(4) => 
                           del_reg_wb_1_4_port, d(3) => del_reg_wb_1_3_port, 
                           d(2) => del_reg_wb_1_2_port, d(1) => 
                           del_reg_wb_1_1_port, d(0) => del_reg_wb_1_0_port, 
                           Q(4) => del_reg_wb_2_4_port, Q(3) => 
                           del_reg_wb_2_3_port, Q(2) => del_reg_wb_2_2_port, 
                           Q(1) => del_reg_wb_2_1_port, Q(0) => 
                           del_reg_wb_2_0_port);
   delay_reg_wb_3 : reg_nbit_n5_1 port map( clk => n2, reset => n1, d(4) => 
                           del_reg_wb_2_4_port, d(3) => del_reg_wb_2_3_port, 
                           d(2) => del_reg_wb_2_2_port, d(1) => 
                           del_reg_wb_2_1_port, d(0) => del_reg_wb_2_0_port, 
                           Q(4) => address_rf_write_4_port, Q(3) => 
                           address_rf_write_3_port, Q(2) => 
                           address_rf_write_2_port, Q(1) => 
                           address_rf_write_1_port, Q(0) => 
                           address_rf_write_0_port);
   reg_file : register_file_NBITREG32_NBITADD5 port map( CLK => n2, RESET => n1
                           , ENABLE => enable_rf_i, RD1 => read_rf_p1, RD2 => 
                           read_rf_p2, WR => write_rf, ADD_WR(4) => 
                           address_rf_write_4_port, ADD_WR(3) => 
                           address_rf_write_3_port, ADD_WR(2) => 
                           address_rf_write_2_port, ADD_WR(1) => 
                           address_rf_write_1_port, ADD_WR(0) => 
                           address_rf_write_0_port, ADD_RD1(4) => 
                           instruction_reg(25), ADD_RD1(3) => 
                           instruction_reg(24), ADD_RD1(2) => 
                           instruction_reg(23), ADD_RD1(1) => 
                           instruction_reg(22), ADD_RD1(0) => 
                           instruction_reg(21), ADD_RD2(4) => 
                           instruction_reg(20), ADD_RD2(3) => 
                           instruction_reg(19), ADD_RD2(2) => 
                           instruction_reg(18), ADD_RD2(1) => 
                           instruction_reg(17), ADD_RD2(0) => 
                           instruction_reg(16), DATAIN(31) => n12, DATAIN(30) 
                           => n13, DATAIN(29) => n14, DATAIN(28) => n15, 
                           DATAIN(27) => n16, DATAIN(26) => n17, DATAIN(25) => 
                           n18, DATAIN(24) => n19, DATAIN(23) => n20, 
                           DATAIN(22) => n21, DATAIN(21) => n22, DATAIN(20) => 
                           n23, DATAIN(19) => n24, DATAIN(18) => n25, 
                           DATAIN(17) => n26, DATAIN(16) => n27, DATAIN(15) => 
                           n28, DATAIN(14) => n29, DATAIN(13) => n30, 
                           DATAIN(12) => n31, DATAIN(11) => n32, DATAIN(10) => 
                           n33, DATAIN(9) => n34, DATAIN(8) => n35, DATAIN(7) 
                           => n36, DATAIN(6) => n37, DATAIN(5) => n38, 
                           DATAIN(4) => n39, DATAIN(3) => n40, DATAIN(2) => n41
                           , DATAIN(1) => n42, DATAIN(0) => n43, OUT1(31) => 
                           val_reg_a_i_31_port, OUT1(30) => val_reg_a_i_30_port
                           , OUT1(29) => val_reg_a_i_29_port, OUT1(28) => 
                           val_reg_a_i_28_port, OUT1(27) => val_reg_a_i_27_port
                           , OUT1(26) => val_reg_a_i_26_port, OUT1(25) => 
                           val_reg_a_i_25_port, OUT1(24) => val_reg_a_i_24_port
                           , OUT1(23) => val_reg_a_i_23_port, OUT1(22) => 
                           val_reg_a_i_22_port, OUT1(21) => val_reg_a_i_21_port
                           , OUT1(20) => val_reg_a_i_20_port, OUT1(19) => 
                           val_reg_a_i_19_port, OUT1(18) => val_reg_a_i_18_port
                           , OUT1(17) => val_reg_a_i_17_port, OUT1(16) => 
                           val_reg_a_i_16_port, OUT1(15) => val_reg_a_i_15_port
                           , OUT1(14) => val_reg_a_i_14_port, OUT1(13) => 
                           val_reg_a_i_13_port, OUT1(12) => val_reg_a_i_12_port
                           , OUT1(11) => val_reg_a_i_11_port, OUT1(10) => 
                           val_reg_a_i_10_port, OUT1(9) => val_reg_a_i_9_port, 
                           OUT1(8) => val_reg_a_i_8_port, OUT1(7) => 
                           val_reg_a_i_7_port, OUT1(6) => val_reg_a_i_6_port, 
                           OUT1(5) => val_reg_a_i_5_port, OUT1(4) => 
                           val_reg_a_i_4_port, OUT1(3) => val_reg_a_i_3_port, 
                           OUT1(2) => val_reg_a_i_2_port, OUT1(1) => 
                           val_reg_a_i_1_port, OUT1(0) => val_reg_a_i_0_port, 
                           OUT2(31) => val_reg_b_i_31_port, OUT2(30) => 
                           val_reg_b_i_30_port, OUT2(29) => val_reg_b_i_29_port
                           , OUT2(28) => val_reg_b_i_28_port, OUT2(27) => 
                           val_reg_b_i_27_port, OUT2(26) => val_reg_b_i_26_port
                           , OUT2(25) => val_reg_b_i_25_port, OUT2(24) => 
                           val_reg_b_i_24_port, OUT2(23) => val_reg_b_i_23_port
                           , OUT2(22) => val_reg_b_i_22_port, OUT2(21) => 
                           val_reg_b_i_21_port, OUT2(20) => val_reg_b_i_20_port
                           , OUT2(19) => val_reg_b_i_19_port, OUT2(18) => 
                           val_reg_b_i_18_port, OUT2(17) => val_reg_b_i_17_port
                           , OUT2(16) => val_reg_b_i_16_port, OUT2(15) => 
                           val_reg_b_i_15_port, OUT2(14) => val_reg_b_i_14_port
                           , OUT2(13) => val_reg_b_i_13_port, OUT2(12) => 
                           val_reg_b_i_12_port, OUT2(11) => val_reg_b_i_11_port
                           , OUT2(10) => val_reg_b_i_10_port, OUT2(9) => 
                           val_reg_b_i_9_port, OUT2(8) => val_reg_b_i_8_port, 
                           OUT2(7) => val_reg_b_i_7_port, OUT2(6) => 
                           val_reg_b_i_6_port, OUT2(5) => val_reg_b_i_5_port, 
                           OUT2(4) => val_reg_b_i_4_port, OUT2(3) => 
                           val_reg_b_i_3_port, OUT2(2) => val_reg_b_i_2_port, 
                           OUT2(1) => val_reg_b_i_1_port, OUT2(0) => 
                           val_reg_b_i_0_port);
   reg_a : reg_nbit_n32_13 port map( clk => n2, reset => n1, d(31) => 
                           val_reg_a_i_31_port, d(30) => val_reg_a_i_30_port, 
                           d(29) => val_reg_a_i_29_port, d(28) => 
                           val_reg_a_i_28_port, d(27) => val_reg_a_i_27_port, 
                           d(26) => val_reg_a_i_26_port, d(25) => 
                           val_reg_a_i_25_port, d(24) => val_reg_a_i_24_port, 
                           d(23) => val_reg_a_i_23_port, d(22) => 
                           val_reg_a_i_22_port, d(21) => val_reg_a_i_21_port, 
                           d(20) => val_reg_a_i_20_port, d(19) => 
                           val_reg_a_i_19_port, d(18) => val_reg_a_i_18_port, 
                           d(17) => val_reg_a_i_17_port, d(16) => 
                           val_reg_a_i_16_port, d(15) => val_reg_a_i_15_port, 
                           d(14) => val_reg_a_i_14_port, d(13) => 
                           val_reg_a_i_13_port, d(12) => val_reg_a_i_12_port, 
                           d(11) => val_reg_a_i_11_port, d(10) => 
                           val_reg_a_i_10_port, d(9) => val_reg_a_i_9_port, 
                           d(8) => val_reg_a_i_8_port, d(7) => 
                           val_reg_a_i_7_port, d(6) => val_reg_a_i_6_port, d(5)
                           => val_reg_a_i_5_port, d(4) => val_reg_a_i_4_port, 
                           d(3) => val_reg_a_i_3_port, d(2) => 
                           val_reg_a_i_2_port, d(1) => val_reg_a_i_1_port, d(0)
                           => val_reg_a_i_0_port, Q(31) => val_a(31), Q(30) => 
                           val_a(30), Q(29) => val_a(29), Q(28) => val_a(28), 
                           Q(27) => val_a(27), Q(26) => val_a(26), Q(25) => 
                           val_a(25), Q(24) => val_a(24), Q(23) => val_a(23), 
                           Q(22) => val_a(22), Q(21) => val_a(21), Q(20) => 
                           val_a(20), Q(19) => val_a(19), Q(18) => val_a(18), 
                           Q(17) => val_a(17), Q(16) => val_a(16), Q(15) => 
                           val_a(15), Q(14) => val_a(14), Q(13) => val_a(13), 
                           Q(12) => val_a(12), Q(11) => val_a(11), Q(10) => 
                           val_a(10), Q(9) => val_a(9), Q(8) => val_a(8), Q(7) 
                           => val_a(7), Q(6) => val_a(6), Q(5) => val_a(5), 
                           Q(4) => val_a(4), Q(3) => val_a(3), Q(2) => val_a(2)
                           , Q(1) => val_a(1), Q(0) => val_a(0));
   reg_b : reg_nbit_n32_12 port map( clk => n2, reset => n1, d(31) => 
                           val_reg_b_i_31_port, d(30) => val_reg_b_i_30_port, 
                           d(29) => val_reg_b_i_29_port, d(28) => 
                           val_reg_b_i_28_port, d(27) => val_reg_b_i_27_port, 
                           d(26) => val_reg_b_i_26_port, d(25) => 
                           val_reg_b_i_25_port, d(24) => val_reg_b_i_24_port, 
                           d(23) => val_reg_b_i_23_port, d(22) => 
                           val_reg_b_i_22_port, d(21) => val_reg_b_i_21_port, 
                           d(20) => val_reg_b_i_20_port, d(19) => 
                           val_reg_b_i_19_port, d(18) => val_reg_b_i_18_port, 
                           d(17) => val_reg_b_i_17_port, d(16) => 
                           val_reg_b_i_16_port, d(15) => val_reg_b_i_15_port, 
                           d(14) => val_reg_b_i_14_port, d(13) => 
                           val_reg_b_i_13_port, d(12) => val_reg_b_i_12_port, 
                           d(11) => val_reg_b_i_11_port, d(10) => 
                           val_reg_b_i_10_port, d(9) => val_reg_b_i_9_port, 
                           d(8) => val_reg_b_i_8_port, d(7) => 
                           val_reg_b_i_7_port, d(6) => val_reg_b_i_6_port, d(5)
                           => val_reg_b_i_5_port, d(4) => val_reg_b_i_4_port, 
                           d(3) => val_reg_b_i_3_port, d(2) => 
                           val_reg_b_i_2_port, d(1) => val_reg_b_i_1_port, d(0)
                           => val_reg_b_i_0_port, Q(31) => val_b(31), Q(30) => 
                           val_b(30), Q(29) => val_b(29), Q(28) => val_b(28), 
                           Q(27) => val_b(27), Q(26) => val_b(26), Q(25) => 
                           val_b(25), Q(24) => val_b(24), Q(23) => val_b(23), 
                           Q(22) => val_b(22), Q(21) => val_b(21), Q(20) => 
                           val_b(20), Q(19) => val_b(19), Q(18) => val_b(18), 
                           Q(17) => val_b(17), Q(16) => val_b(16), Q(15) => 
                           val_b(15), Q(14) => val_b(14), Q(13) => val_b(13), 
                           Q(12) => val_b(12), Q(11) => val_b(11), Q(10) => 
                           val_b(10), Q(9) => val_b(9), Q(8) => val_b(8), Q(7) 
                           => val_b(7), Q(6) => val_b(6), Q(5) => val_b(5), 
                           Q(4) => val_b(4), Q(3) => val_b(3), Q(2) => val_b(2)
                           , Q(1) => val_b(1), Q(0) => val_b(0));
   sign_extension_logic_immediate : sign_extension_N32_STARTING_BIT16 port map(
                           val_to_exetend(15) => instruction_reg(15), 
                           val_to_exetend(14) => instruction_reg(14), 
                           val_to_exetend(13) => instruction_reg(13), 
                           val_to_exetend(12) => instruction_reg(12), 
                           val_to_exetend(11) => instruction_reg(11), 
                           val_to_exetend(10) => instruction_reg(10), 
                           val_to_exetend(9) => instruction_reg(9), 
                           val_to_exetend(8) => instruction_reg(8), 
                           val_to_exetend(7) => instruction_reg(7), 
                           val_to_exetend(6) => instruction_reg(6), 
                           val_to_exetend(5) => instruction_reg(5), 
                           val_to_exetend(4) => instruction_reg(4), 
                           val_to_exetend(3) => instruction_reg(3), 
                           val_to_exetend(2) => instruction_reg(2), 
                           val_to_exetend(1) => instruction_reg(1), 
                           val_to_exetend(0) => instruction_reg(0), enable => 
                           compute_sext, extended_val(31) => 
                           val_reg_immediate_i_31_port, extended_val(30) => 
                           val_reg_immediate_i_30_port, extended_val(29) => 
                           val_reg_immediate_i_29_port, extended_val(28) => 
                           val_reg_immediate_i_28_port, extended_val(27) => 
                           val_reg_immediate_i_27_port, extended_val(26) => 
                           val_reg_immediate_i_26_port, extended_val(25) => 
                           val_reg_immediate_i_25_port, extended_val(24) => 
                           val_reg_immediate_i_24_port, extended_val(23) => 
                           val_reg_immediate_i_23_port, extended_val(22) => 
                           val_reg_immediate_i_22_port, extended_val(21) => 
                           val_reg_immediate_i_21_port, extended_val(20) => 
                           val_reg_immediate_i_20_port, extended_val(19) => 
                           val_reg_immediate_i_19_port, extended_val(18) => 
                           val_reg_immediate_i_18_port, extended_val(17) => 
                           val_reg_immediate_i_17_port, extended_val(16) => 
                           val_reg_immediate_i_16_port, extended_val(15) => 
                           val_reg_immediate_i_15_port, extended_val(14) => 
                           val_reg_immediate_i_14_port, extended_val(13) => 
                           val_reg_immediate_i_13_port, extended_val(12) => 
                           val_reg_immediate_i_12_port, extended_val(11) => 
                           val_reg_immediate_i_11_port, extended_val(10) => 
                           val_reg_immediate_i_10_port, extended_val(9) => 
                           val_reg_immediate_i_9_port, extended_val(8) => 
                           val_reg_immediate_i_8_port, extended_val(7) => 
                           val_reg_immediate_i_7_port, extended_val(6) => 
                           val_reg_immediate_i_6_port, extended_val(5) => 
                           val_reg_immediate_i_5_port, extended_val(4) => 
                           val_reg_immediate_i_4_port, extended_val(3) => 
                           val_reg_immediate_i_3_port, extended_val(2) => 
                           val_reg_immediate_i_2_port, extended_val(1) => 
                           val_reg_immediate_i_1_port, extended_val(0) => 
                           val_reg_immediate_i_0_port);
   sign_extension_logic_jump : sign_extension_N32_STARTING_BIT26 port map( 
                           val_to_exetend(25) => instruction_reg(25), 
                           val_to_exetend(24) => instruction_reg(24), 
                           val_to_exetend(23) => instruction_reg(23), 
                           val_to_exetend(22) => instruction_reg(22), 
                           val_to_exetend(21) => instruction_reg(21), 
                           val_to_exetend(20) => instruction_reg(20), 
                           val_to_exetend(19) => instruction_reg(19), 
                           val_to_exetend(18) => instruction_reg(18), 
                           val_to_exetend(17) => instruction_reg(17), 
                           val_to_exetend(16) => instruction_reg(16), 
                           val_to_exetend(15) => instruction_reg(15), 
                           val_to_exetend(14) => instruction_reg(14), 
                           val_to_exetend(13) => instruction_reg(13), 
                           val_to_exetend(12) => instruction_reg(12), 
                           val_to_exetend(11) => instruction_reg(11), 
                           val_to_exetend(10) => instruction_reg(10), 
                           val_to_exetend(9) => instruction_reg(9), 
                           val_to_exetend(8) => instruction_reg(8), 
                           val_to_exetend(7) => instruction_reg(7), 
                           val_to_exetend(6) => instruction_reg(6), 
                           val_to_exetend(5) => instruction_reg(5), 
                           val_to_exetend(4) => instruction_reg(4), 
                           val_to_exetend(3) => instruction_reg(3), 
                           val_to_exetend(2) => instruction_reg(2), 
                           val_to_exetend(1) => instruction_reg(1), 
                           val_to_exetend(0) => instruction_reg(0), enable => 
                           enable_sign_extension_logic, extended_val(31) => 
                           val_reg_immediate_j_31_port, extended_val(30) => 
                           val_reg_immediate_j_30_port, extended_val(29) => 
                           val_reg_immediate_j_29_port, extended_val(28) => 
                           val_reg_immediate_j_28_port, extended_val(27) => 
                           val_reg_immediate_j_27_port, extended_val(26) => 
                           val_reg_immediate_j_26_port, extended_val(25) => 
                           val_reg_immediate_j_25_port, extended_val(24) => 
                           val_reg_immediate_j_24_port, extended_val(23) => 
                           val_reg_immediate_j_23_port, extended_val(22) => 
                           val_reg_immediate_j_22_port, extended_val(21) => 
                           val_reg_immediate_j_21_port, extended_val(20) => 
                           val_reg_immediate_j_20_port, extended_val(19) => 
                           val_reg_immediate_j_19_port, extended_val(18) => 
                           val_reg_immediate_j_18_port, extended_val(17) => 
                           val_reg_immediate_j_17_port, extended_val(16) => 
                           val_reg_immediate_j_16_port, extended_val(15) => 
                           val_reg_immediate_j_15_port, extended_val(14) => 
                           val_reg_immediate_j_14_port, extended_val(13) => 
                           val_reg_immediate_j_13_port, extended_val(12) => 
                           val_reg_immediate_j_12_port, extended_val(11) => 
                           val_reg_immediate_j_11_port, extended_val(10) => 
                           val_reg_immediate_j_10_port, extended_val(9) => 
                           val_reg_immediate_j_9_port, extended_val(8) => 
                           val_reg_immediate_j_8_port, extended_val(7) => 
                           val_reg_immediate_j_7_port, extended_val(6) => 
                           val_reg_immediate_j_6_port, extended_val(5) => 
                           val_reg_immediate_j_5_port, extended_val(4) => 
                           val_reg_immediate_j_4_port, extended_val(3) => 
                           val_reg_immediate_j_3_port, extended_val(2) => 
                           val_reg_immediate_j_2_port, extended_val(1) => 
                           val_reg_immediate_j_1_port, extended_val(0) => 
                           val_reg_immediate_j_0_port);
   immediate_reg_mux : MUX_zbit_nbit_N32_Z1_0 port map( inputs(0) => 
                           val_reg_immediate_i_31_port, inputs(1) => 
                           val_reg_immediate_i_30_port, inputs(2) => 
                           val_reg_immediate_i_29_port, inputs(3) => 
                           val_reg_immediate_i_28_port, inputs(4) => 
                           val_reg_immediate_i_27_port, inputs(5) => 
                           val_reg_immediate_i_26_port, inputs(6) => 
                           val_reg_immediate_i_25_port, inputs(7) => 
                           val_reg_immediate_i_24_port, inputs(8) => 
                           val_reg_immediate_i_23_port, inputs(9) => 
                           val_reg_immediate_i_22_port, inputs(10) => 
                           val_reg_immediate_i_21_port, inputs(11) => 
                           val_reg_immediate_i_20_port, inputs(12) => 
                           val_reg_immediate_i_19_port, inputs(13) => 
                           val_reg_immediate_i_18_port, inputs(14) => 
                           val_reg_immediate_i_17_port, inputs(15) => 
                           val_reg_immediate_i_16_port, inputs(16) => 
                           val_reg_immediate_i_15_port, inputs(17) => 
                           val_reg_immediate_i_14_port, inputs(18) => 
                           val_reg_immediate_i_13_port, inputs(19) => 
                           val_reg_immediate_i_12_port, inputs(20) => 
                           val_reg_immediate_i_11_port, inputs(21) => 
                           val_reg_immediate_i_10_port, inputs(22) => 
                           val_reg_immediate_i_9_port, inputs(23) => 
                           val_reg_immediate_i_8_port, inputs(24) => 
                           val_reg_immediate_i_7_port, inputs(25) => 
                           val_reg_immediate_i_6_port, inputs(26) => 
                           val_reg_immediate_i_5_port, inputs(27) => 
                           val_reg_immediate_i_4_port, inputs(28) => 
                           val_reg_immediate_i_3_port, inputs(29) => 
                           val_reg_immediate_i_2_port, inputs(30) => 
                           val_reg_immediate_i_1_port, inputs(31) => 
                           val_reg_immediate_i_0_port, inputs(32) => 
                           val_reg_immediate_j_31_port, inputs(33) => 
                           val_reg_immediate_j_30_port, inputs(34) => 
                           val_reg_immediate_j_29_port, inputs(35) => 
                           val_reg_immediate_j_28_port, inputs(36) => 
                           val_reg_immediate_j_27_port, inputs(37) => 
                           val_reg_immediate_j_26_port, inputs(38) => 
                           val_reg_immediate_j_25_port, inputs(39) => 
                           val_reg_immediate_j_24_port, inputs(40) => 
                           val_reg_immediate_j_23_port, inputs(41) => 
                           val_reg_immediate_j_22_port, inputs(42) => 
                           val_reg_immediate_j_21_port, inputs(43) => 
                           val_reg_immediate_j_20_port, inputs(44) => 
                           val_reg_immediate_j_19_port, inputs(45) => 
                           val_reg_immediate_j_18_port, inputs(46) => 
                           val_reg_immediate_j_17_port, inputs(47) => 
                           val_reg_immediate_j_16_port, inputs(48) => 
                           val_reg_immediate_j_15_port, inputs(49) => 
                           val_reg_immediate_j_14_port, inputs(50) => 
                           val_reg_immediate_j_13_port, inputs(51) => 
                           val_reg_immediate_j_12_port, inputs(52) => 
                           val_reg_immediate_j_11_port, inputs(53) => 
                           val_reg_immediate_j_10_port, inputs(54) => 
                           val_reg_immediate_j_9_port, inputs(55) => 
                           val_reg_immediate_j_8_port, inputs(56) => 
                           val_reg_immediate_j_7_port, inputs(57) => 
                           val_reg_immediate_j_6_port, inputs(58) => 
                           val_reg_immediate_j_5_port, inputs(59) => 
                           val_reg_immediate_j_4_port, inputs(60) => 
                           val_reg_immediate_j_3_port, inputs(61) => 
                           val_reg_immediate_j_2_port, inputs(62) => 
                           val_reg_immediate_j_1_port, inputs(63) => 
                           val_reg_immediate_j_0_port, SEL => n81, Y(31) => 
                           val_reg_immediate_31_port, Y(30) => 
                           val_reg_immediate_30_port, Y(29) => 
                           val_reg_immediate_29_port, Y(28) => 
                           val_reg_immediate_28_port, Y(27) => 
                           val_reg_immediate_27_port, Y(26) => 
                           val_reg_immediate_26_port, Y(25) => 
                           val_reg_immediate_25_port, Y(24) => 
                           val_reg_immediate_24_port, Y(23) => 
                           val_reg_immediate_23_port, Y(22) => 
                           val_reg_immediate_22_port, Y(21) => 
                           val_reg_immediate_21_port, Y(20) => 
                           val_reg_immediate_20_port, Y(19) => 
                           val_reg_immediate_19_port, Y(18) => 
                           val_reg_immediate_18_port, Y(17) => 
                           val_reg_immediate_17_port, Y(16) => 
                           val_reg_immediate_16_port, Y(15) => 
                           val_reg_immediate_15_port, Y(14) => 
                           val_reg_immediate_14_port, Y(13) => 
                           val_reg_immediate_13_port, Y(12) => 
                           val_reg_immediate_12_port, Y(11) => 
                           val_reg_immediate_11_port, Y(10) => 
                           val_reg_immediate_10_port, Y(9) => 
                           val_reg_immediate_9_port, Y(8) => 
                           val_reg_immediate_8_port, Y(7) => 
                           val_reg_immediate_7_port, Y(6) => 
                           val_reg_immediate_6_port, Y(5) => 
                           val_reg_immediate_5_port, Y(4) => 
                           val_reg_immediate_4_port, Y(3) => 
                           val_reg_immediate_3_port, Y(2) => 
                           val_reg_immediate_2_port, Y(1) => 
                           val_reg_immediate_1_port, Y(0) => 
                           val_reg_immediate_0_port);
   reg_immediate : reg_nbit_n32_11 port map( clk => clk_immediate, reset => n1,
                           d(31) => val_reg_immediate_31_port, d(30) => 
                           val_reg_immediate_30_port, d(29) => 
                           val_reg_immediate_29_port, d(28) => 
                           val_reg_immediate_28_port, d(27) => 
                           val_reg_immediate_27_port, d(26) => 
                           val_reg_immediate_26_port, d(25) => 
                           val_reg_immediate_25_port, d(24) => 
                           val_reg_immediate_24_port, d(23) => 
                           val_reg_immediate_23_port, d(22) => 
                           val_reg_immediate_22_port, d(21) => 
                           val_reg_immediate_21_port, d(20) => 
                           val_reg_immediate_20_port, d(19) => 
                           val_reg_immediate_19_port, d(18) => 
                           val_reg_immediate_18_port, d(17) => 
                           val_reg_immediate_17_port, d(16) => 
                           val_reg_immediate_16_port, d(15) => 
                           val_reg_immediate_15_port, d(14) => 
                           val_reg_immediate_14_port, d(13) => 
                           val_reg_immediate_13_port, d(12) => 
                           val_reg_immediate_12_port, d(11) => 
                           val_reg_immediate_11_port, d(10) => 
                           val_reg_immediate_10_port, d(9) => 
                           val_reg_immediate_9_port, d(8) => 
                           val_reg_immediate_8_port, d(7) => 
                           val_reg_immediate_7_port, d(6) => 
                           val_reg_immediate_6_port, d(5) => 
                           val_reg_immediate_5_port, d(4) => 
                           val_reg_immediate_4_port, d(3) => 
                           val_reg_immediate_3_port, d(2) => 
                           val_reg_immediate_2_port, d(1) => 
                           val_reg_immediate_1_port, d(0) => 
                           val_reg_immediate_0_port, Q(31) => val_immediate(31)
                           , Q(30) => val_immediate(30), Q(29) => 
                           val_immediate(29), Q(28) => val_immediate(28), Q(27)
                           => val_immediate(27), Q(26) => val_immediate(26), 
                           Q(25) => val_immediate(25), Q(24) => 
                           val_immediate(24), Q(23) => val_immediate(23), Q(22)
                           => val_immediate(22), Q(21) => val_immediate(21), 
                           Q(20) => val_immediate(20), Q(19) => 
                           val_immediate(19), Q(18) => val_immediate(18), Q(17)
                           => val_immediate(17), Q(16) => val_immediate(16), 
                           Q(15) => val_immediate(15), Q(14) => 
                           val_immediate(14), Q(13) => val_immediate(13), Q(12)
                           => val_immediate(12), Q(11) => val_immediate(11), 
                           Q(10) => val_immediate(10), Q(9) => val_immediate(9)
                           , Q(8) => val_immediate(8), Q(7) => val_immediate(7)
                           , Q(6) => val_immediate(6), Q(5) => val_immediate(5)
                           , Q(4) => val_immediate(4), Q(3) => val_immediate(3)
                           , Q(2) => val_immediate(2), Q(1) => val_immediate(1)
                           , Q(0) => val_immediate(0));
   pc_delay_reg1 : reg_nbit_n33_0 port map( clk => n2, reset => n1, d(32) => 
                           new_prog_counter_val(31), d(31) => 
                           new_prog_counter_val(30), d(30) => 
                           new_prog_counter_val(29), d(29) => 
                           new_prog_counter_val(28), d(28) => 
                           new_prog_counter_val(27), d(27) => 
                           new_prog_counter_val(26), d(26) => 
                           new_prog_counter_val(25), d(25) => 
                           new_prog_counter_val(24), d(24) => 
                           new_prog_counter_val(23), d(23) => 
                           new_prog_counter_val(22), d(22) => 
                           new_prog_counter_val(21), d(21) => 
                           new_prog_counter_val(20), d(20) => 
                           new_prog_counter_val(19), d(19) => 
                           new_prog_counter_val(18), d(18) => 
                           new_prog_counter_val(17), d(17) => 
                           new_prog_counter_val(16), d(16) => 
                           new_prog_counter_val(15), d(15) => 
                           new_prog_counter_val(14), d(14) => 
                           new_prog_counter_val(13), d(13) => 
                           new_prog_counter_val(12), d(12) => 
                           new_prog_counter_val(11), d(11) => 
                           new_prog_counter_val(10), d(10) => 
                           new_prog_counter_val(9), d(9) => 
                           new_prog_counter_val(8), d(8) => 
                           new_prog_counter_val(7), d(7) => 
                           new_prog_counter_val(6), d(6) => 
                           new_prog_counter_val(5), d(5) => 
                           new_prog_counter_val(4), d(4) => 
                           new_prog_counter_val(3), d(3) => 
                           new_prog_counter_val(2), d(2) => 
                           new_prog_counter_val(1), d(1) => 
                           new_prog_counter_val(0), d(0) => jump_sext, Q(32) =>
                           pc_delay2_32_port, Q(31) => pc_delay2_31_port, Q(30)
                           => pc_delay2_30_port, Q(29) => pc_delay2_29_port, 
                           Q(28) => pc_delay2_28_port, Q(27) => 
                           pc_delay2_27_port, Q(26) => pc_delay2_26_port, Q(25)
                           => pc_delay2_25_port, Q(24) => pc_delay2_24_port, 
                           Q(23) => pc_delay2_23_port, Q(22) => 
                           pc_delay2_22_port, Q(21) => pc_delay2_21_port, Q(20)
                           => pc_delay2_20_port, Q(19) => pc_delay2_19_port, 
                           Q(18) => pc_delay2_18_port, Q(17) => 
                           pc_delay2_17_port, Q(16) => pc_delay2_16_port, Q(15)
                           => pc_delay2_15_port, Q(14) => pc_delay2_14_port, 
                           Q(13) => pc_delay2_13_port, Q(12) => 
                           pc_delay2_12_port, Q(11) => pc_delay2_11_port, Q(10)
                           => pc_delay2_10_port, Q(9) => pc_delay2_9_port, Q(8)
                           => pc_delay2_8_port, Q(7) => pc_delay2_7_port, Q(6) 
                           => pc_delay2_6_port, Q(5) => pc_delay2_5_port, Q(4) 
                           => pc_delay2_4_port, Q(3) => pc_delay2_3_port, Q(2) 
                           => pc_delay2_2_port, Q(1) => pc_delay2_1_port, Q(0) 
                           => pc_delay2_0_port);
   pc_delay_reg_2 : reg_nbit_n33_1 port map( clk => n2, reset => n1, d(32) => 
                           pc_delay2_32_port, d(31) => pc_delay2_31_port, d(30)
                           => pc_delay2_30_port, d(29) => pc_delay2_29_port, 
                           d(28) => pc_delay2_28_port, d(27) => 
                           pc_delay2_27_port, d(26) => pc_delay2_26_port, d(25)
                           => pc_delay2_25_port, d(24) => pc_delay2_24_port, 
                           d(23) => pc_delay2_23_port, d(22) => 
                           pc_delay2_22_port, d(21) => pc_delay2_21_port, d(20)
                           => pc_delay2_20_port, d(19) => pc_delay2_19_port, 
                           d(18) => pc_delay2_18_port, d(17) => 
                           pc_delay2_17_port, d(16) => pc_delay2_16_port, d(15)
                           => pc_delay2_15_port, d(14) => pc_delay2_14_port, 
                           d(13) => pc_delay2_13_port, d(12) => 
                           pc_delay2_12_port, d(11) => pc_delay2_11_port, d(10)
                           => pc_delay2_10_port, d(9) => pc_delay2_9_port, d(8)
                           => pc_delay2_8_port, d(7) => pc_delay2_7_port, d(6) 
                           => pc_delay2_6_port, d(5) => pc_delay2_5_port, d(4) 
                           => pc_delay2_4_port, d(3) => pc_delay2_3_port, d(2) 
                           => pc_delay2_2_port, d(1) => pc_delay2_1_port, d(0) 
                           => pc_delay2_0_port, Q(32) => pc_delay3_32_port, 
                           Q(31) => pc_delay3_31_port, Q(30) => 
                           pc_delay3_30_port, Q(29) => pc_delay3_29_port, Q(28)
                           => pc_delay3_28_port, Q(27) => pc_delay3_27_port, 
                           Q(26) => pc_delay3_26_port, Q(25) => 
                           pc_delay3_25_port, Q(24) => pc_delay3_24_port, Q(23)
                           => pc_delay3_23_port, Q(22) => pc_delay3_22_port, 
                           Q(21) => pc_delay3_21_port, Q(20) => 
                           pc_delay3_20_port, Q(19) => pc_delay3_19_port, Q(18)
                           => pc_delay3_18_port, Q(17) => pc_delay3_17_port, 
                           Q(16) => pc_delay3_16_port, Q(15) => 
                           pc_delay3_15_port, Q(14) => pc_delay3_14_port, Q(13)
                           => pc_delay3_13_port, Q(12) => pc_delay3_12_port, 
                           Q(11) => pc_delay3_11_port, Q(10) => 
                           pc_delay3_10_port, Q(9) => pc_delay3_9_port, Q(8) =>
                           pc_delay3_8_port, Q(7) => pc_delay3_7_port, Q(6) => 
                           pc_delay3_6_port, Q(5) => pc_delay3_5_port, Q(4) => 
                           pc_delay3_4_port, Q(3) => pc_delay3_3_port, Q(2) => 
                           pc_delay3_2_port, Q(1) => pc_delay3_1_port, Q(0) => 
                           pc_delay3_0_port);
   U2 : AND3_X2 port map( A1 => address_rf_write_4_port, A2 => 
                           address_rf_write_3_port, A3 => n4, ZN => n3);
   U3 : INV_X2 port map( A => compute_sext, ZN => n81);
   U4 : AOI211_X4 port map( C1 => n10, C2 => enable_rf, A => n81, B => n11, ZN 
                           => enable_sign_extension_logic);
   U5 : BUF_X2 port map( A => n82, Z => n1);
   U6 : BUF_X1 port map( A => clk, Z => n2);
   U7 : MUX2_X1 port map( A => update_reg_value(31), B => pc_delay3_32_port, S 
                           => n3, Z => n12);
   U8 : MUX2_X1 port map( A => update_reg_value(30), B => pc_delay3_31_port, S 
                           => n3, Z => n13);
   U9 : MUX2_X1 port map( A => update_reg_value(29), B => pc_delay3_30_port, S 
                           => n3, Z => n14);
   U10 : MUX2_X1 port map( A => update_reg_value(28), B => pc_delay3_29_port, S
                           => n3, Z => n15);
   U11 : MUX2_X1 port map( A => update_reg_value(27), B => pc_delay3_28_port, S
                           => n3, Z => n16);
   U12 : MUX2_X1 port map( A => update_reg_value(26), B => pc_delay3_27_port, S
                           => n3, Z => n17);
   U13 : MUX2_X1 port map( A => update_reg_value(25), B => pc_delay3_26_port, S
                           => n3, Z => n18);
   U14 : MUX2_X1 port map( A => update_reg_value(24), B => pc_delay3_25_port, S
                           => n3, Z => n19);
   U15 : MUX2_X1 port map( A => update_reg_value(23), B => pc_delay3_24_port, S
                           => n3, Z => n20);
   U16 : MUX2_X1 port map( A => update_reg_value(22), B => pc_delay3_23_port, S
                           => n3, Z => n21);
   U17 : MUX2_X1 port map( A => update_reg_value(21), B => pc_delay3_22_port, S
                           => n3, Z => n22);
   U18 : MUX2_X1 port map( A => update_reg_value(20), B => pc_delay3_21_port, S
                           => n3, Z => n23);
   U19 : MUX2_X1 port map( A => update_reg_value(19), B => pc_delay3_20_port, S
                           => n3, Z => n24);
   U20 : MUX2_X1 port map( A => update_reg_value(18), B => pc_delay3_19_port, S
                           => n3, Z => n25);
   U21 : MUX2_X1 port map( A => update_reg_value(17), B => pc_delay3_18_port, S
                           => n3, Z => n26);
   U22 : MUX2_X1 port map( A => update_reg_value(16), B => pc_delay3_17_port, S
                           => n3, Z => n27);
   U23 : MUX2_X1 port map( A => update_reg_value(15), B => pc_delay3_16_port, S
                           => n3, Z => n28);
   U24 : MUX2_X1 port map( A => update_reg_value(14), B => pc_delay3_15_port, S
                           => n3, Z => n29);
   U25 : MUX2_X1 port map( A => update_reg_value(13), B => pc_delay3_14_port, S
                           => n3, Z => n30);
   U26 : MUX2_X1 port map( A => update_reg_value(12), B => pc_delay3_13_port, S
                           => n3, Z => n31);
   U27 : MUX2_X1 port map( A => update_reg_value(11), B => pc_delay3_12_port, S
                           => n3, Z => n32);
   U28 : MUX2_X1 port map( A => update_reg_value(10), B => pc_delay3_11_port, S
                           => n3, Z => n33);
   U29 : MUX2_X1 port map( A => update_reg_value(9), B => pc_delay3_10_port, S 
                           => n3, Z => n34);
   U30 : MUX2_X1 port map( A => update_reg_value(8), B => pc_delay3_9_port, S 
                           => n3, Z => n35);
   U31 : MUX2_X1 port map( A => update_reg_value(7), B => pc_delay3_8_port, S 
                           => n3, Z => n36);
   U32 : MUX2_X1 port map( A => update_reg_value(6), B => pc_delay3_7_port, S 
                           => n3, Z => n37);
   U33 : MUX2_X1 port map( A => update_reg_value(5), B => pc_delay3_6_port, S 
                           => n3, Z => n38);
   U34 : MUX2_X1 port map( A => update_reg_value(4), B => pc_delay3_5_port, S 
                           => n3, Z => n39);
   U35 : MUX2_X1 port map( A => update_reg_value(3), B => pc_delay3_4_port, S 
                           => n3, Z => n40);
   U36 : MUX2_X1 port map( A => update_reg_value(2), B => pc_delay3_3_port, S 
                           => n3, Z => n41);
   U37 : MUX2_X1 port map( A => update_reg_value(1), B => pc_delay3_2_port, S 
                           => n3, Z => n42);
   U38 : MUX2_X1 port map( A => update_reg_value(0), B => pc_delay3_1_port, S 
                           => n3, Z => n43);
   U39 : AND3_X1 port map( A1 => address_rf_write_1_port, A2 => 
                           address_rf_write_0_port, A3 => 
                           address_rf_write_2_port, ZN => n4);
   U40 : MUX2_X1 port map( A => new_prog_counter_val(0), B => pc_delay3_1_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(0));
   U41 : MUX2_X1 port map( A => new_prog_counter_val(1), B => pc_delay3_2_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(1));
   U42 : MUX2_X1 port map( A => new_prog_counter_val(2), B => pc_delay3_3_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(2));
   U43 : MUX2_X1 port map( A => new_prog_counter_val(3), B => pc_delay3_4_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(3));
   U44 : MUX2_X1 port map( A => new_prog_counter_val(4), B => pc_delay3_5_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(4));
   U45 : MUX2_X1 port map( A => new_prog_counter_val(5), B => pc_delay3_6_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(5));
   U46 : MUX2_X1 port map( A => new_prog_counter_val(6), B => pc_delay3_7_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(6));
   U47 : MUX2_X1 port map( A => new_prog_counter_val(7), B => pc_delay3_8_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(7));
   U48 : MUX2_X1 port map( A => new_prog_counter_val(8), B => pc_delay3_9_port,
                           S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(8));
   U49 : MUX2_X1 port map( A => new_prog_counter_val(9), B => pc_delay3_10_port
                           , S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(9));
   U50 : MUX2_X1 port map( A => new_prog_counter_val(10), B => 
                           pc_delay3_11_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(10));
   U51 : MUX2_X1 port map( A => new_prog_counter_val(11), B => 
                           pc_delay3_12_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(11));
   U52 : MUX2_X1 port map( A => new_prog_counter_val(12), B => 
                           pc_delay3_13_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(12));
   U53 : MUX2_X1 port map( A => new_prog_counter_val(13), B => 
                           pc_delay3_14_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(13));
   U54 : MUX2_X1 port map( A => new_prog_counter_val(14), B => 
                           pc_delay3_15_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(14));
   U55 : MUX2_X1 port map( A => new_prog_counter_val(15), B => 
                           pc_delay3_16_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(15));
   U56 : MUX2_X1 port map( A => new_prog_counter_val(16), B => 
                           pc_delay3_17_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(16));
   U57 : MUX2_X1 port map( A => new_prog_counter_val(17), B => 
                           pc_delay3_18_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(17));
   U58 : MUX2_X1 port map( A => new_prog_counter_val(18), B => 
                           pc_delay3_19_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(18));
   U59 : MUX2_X1 port map( A => new_prog_counter_val(19), B => 
                           pc_delay3_20_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(19));
   U60 : MUX2_X1 port map( A => new_prog_counter_val(20), B => 
                           pc_delay3_21_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(20));
   U61 : MUX2_X1 port map( A => new_prog_counter_val(21), B => 
                           pc_delay3_22_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(21));
   U62 : MUX2_X1 port map( A => new_prog_counter_val(22), B => 
                           pc_delay3_23_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(22));
   U63 : MUX2_X1 port map( A => new_prog_counter_val(23), B => 
                           pc_delay3_24_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(23));
   U64 : MUX2_X1 port map( A => new_prog_counter_val(24), B => 
                           pc_delay3_25_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(24));
   U65 : MUX2_X1 port map( A => new_prog_counter_val(25), B => 
                           pc_delay3_26_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(25));
   U66 : MUX2_X1 port map( A => new_prog_counter_val(26), B => 
                           pc_delay3_27_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(26));
   U67 : MUX2_X1 port map( A => new_prog_counter_val(27), B => 
                           pc_delay3_28_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(27));
   U68 : MUX2_X1 port map( A => new_prog_counter_val(28), B => 
                           pc_delay3_29_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(28));
   U69 : MUX2_X1 port map( A => new_prog_counter_val(29), B => 
                           pc_delay3_30_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(29));
   U70 : MUX2_X1 port map( A => new_prog_counter_val(30), B => 
                           pc_delay3_31_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(30));
   U71 : MUX2_X1 port map( A => new_prog_counter_val(31), B => 
                           pc_delay3_32_port, S => pc_delay3_0_port, Z => 
                           new_prog_counter_val_exe(31));
   U72 : OR2_X1 port map( A1 => enable_sign_extension_logic, A2 => n5, ZN => 
                           n76);
   U73 : MUX2_X1 port map( A => instruction_reg(16), B => instruction_reg(11), 
                           S => rtype_itypen, Z => n5);
   U74 : OR2_X1 port map( A1 => enable_sign_extension_logic, A2 => n6, ZN => 
                           n77);
   U75 : MUX2_X1 port map( A => instruction_reg(17), B => instruction_reg(12), 
                           S => rtype_itypen, Z => n6);
   U76 : OR2_X1 port map( A1 => enable_sign_extension_logic, A2 => n7, ZN => 
                           n78);
   U77 : MUX2_X1 port map( A => instruction_reg(18), B => instruction_reg(13), 
                           S => rtype_itypen, Z => n7);
   U78 : OR2_X1 port map( A1 => enable_sign_extension_logic, A2 => n8, ZN => 
                           n79);
   U79 : MUX2_X1 port map( A => instruction_reg(19), B => instruction_reg(14), 
                           S => rtype_itypen, Z => n8);
   U80 : OR2_X1 port map( A1 => enable_sign_extension_logic, A2 => n9, ZN => 
                           n80);
   U81 : MUX2_X1 port map( A => instruction_reg(20), B => instruction_reg(15), 
                           S => rtype_itypen, Z => n9);
   U82 : INV_X1 port map( A => rst, ZN => n82);
   U83 : INV_X1 port map( A => jump_sext, ZN => n11);
   U84 : OR2_X1 port map( A1 => read_rf_p2, A2 => read_rf_p1, ZN => n10);
   U85 : OR2_X1 port map( A1 => enable_rf, A2 => write_rf, ZN => enable_rf_i);
   U86 : AND2_X1 port map( A1 => n2, A2 => compute_sext, ZN => clk_immediate);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity fetch_stage_IR_SIZE32_PC_SIZE32 is

   port( clk, rst : in std_logic;  new_pc_value_mem_stage : in std_logic_vector
         (31 downto 0);  branch_taken : in std_logic;  new_pc_value, 
         IRAM_ADDRESS : out std_logic_vector (31 downto 0);  IRAM_ENABLE : out 
         std_logic;  IRAM_READY : in std_logic;  IRAM_DATA : in 
         std_logic_vector (0 to 31);  curr_instruction : out std_logic_vector 
         (31 downto 0);  iram_enable_cu, update_pc_branch, stall : in std_logic
         ;  iram_ready_cu : out std_logic);

end fetch_stage_IR_SIZE32_PC_SIZE32;

architecture SYN_structural of fetch_stage_IR_SIZE32_PC_SIZE32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component reg_nbit_n32_14
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_15
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_nbit_n32_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (31 downto 0); 
            Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, curr_instruction_31_port, 
      curr_instruction_30_port, curr_instruction_29_port, 
      curr_instruction_28_port, curr_instruction_27_port, 
      curr_instruction_26_port, curr_instruction_25_port, 
      curr_instruction_24_port, curr_instruction_23_port, 
      curr_instruction_22_port, curr_instruction_21_port, 
      curr_instruction_20_port, curr_instruction_19_port, 
      curr_instruction_18_port, curr_instruction_17_port, 
      curr_instruction_16_port, curr_instruction_15_port, 
      curr_instruction_14_port, curr_instruction_13_port, 
      curr_instruction_12_port, curr_instruction_11_port, 
      curr_instruction_10_port, curr_instruction_9_port, 
      curr_instruction_8_port, curr_instruction_7_port, curr_instruction_6_port
      , curr_instruction_5_port, curr_instruction_4_port, 
      curr_instruction_3_port, curr_instruction_2_port, curr_instruction_1_port
      , curr_instruction_0_port, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, 
      N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29
      , N30, N31, N32, N33, N34, N35, N36, N39, N40, N41, N42, N43, N44, N45, 
      N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60
      , N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, n5_port, n6_port, 
      n7_port, n8_port, n1, n2, n3, n4, n9_port, n10_port, n11_port, n12_port, 
      n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, n19_port, 
      n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37, n38, n39_port, n40_port, n41_port, 
      n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, 
      n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, 
      n70_port, n_5534, n_5535 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   IRAM_ENABLE <= iram_enable_cu;
   curr_instruction <= ( curr_instruction_31_port, curr_instruction_30_port, 
      curr_instruction_29_port, curr_instruction_28_port, 
      curr_instruction_27_port, curr_instruction_26_port, 
      curr_instruction_25_port, curr_instruction_24_port, 
      curr_instruction_23_port, curr_instruction_22_port, 
      curr_instruction_21_port, curr_instruction_20_port, 
      curr_instruction_19_port, curr_instruction_18_port, 
      curr_instruction_17_port, curr_instruction_16_port, 
      curr_instruction_15_port, curr_instruction_14_port, 
      curr_instruction_13_port, curr_instruction_12_port, 
      curr_instruction_11_port, curr_instruction_10_port, 
      curr_instruction_9_port, curr_instruction_8_port, curr_instruction_7_port
      , curr_instruction_6_port, curr_instruction_5_port, 
      curr_instruction_4_port, curr_instruction_3_port, curr_instruction_2_port
      , curr_instruction_1_port, curr_instruction_0_port );
   iram_ready_cu <= IRAM_READY;
   
   n5_port <= '0';
   n6_port <= '1';
   n7_port <= '0';
   n8_port <= '0';
   program_counter : reg_nbit_n32_0 port map( clk => clk, reset => n70_port, 
                           d(31) => new_pc_value_mem_stage(31), d(30) => 
                           new_pc_value_mem_stage(30), d(29) => 
                           new_pc_value_mem_stage(29), d(28) => 
                           new_pc_value_mem_stage(28), d(27) => 
                           new_pc_value_mem_stage(27), d(26) => 
                           new_pc_value_mem_stage(26), d(25) => 
                           new_pc_value_mem_stage(25), d(24) => 
                           new_pc_value_mem_stage(24), d(23) => 
                           new_pc_value_mem_stage(23), d(22) => 
                           new_pc_value_mem_stage(22), d(21) => 
                           new_pc_value_mem_stage(21), d(20) => 
                           new_pc_value_mem_stage(20), d(19) => 
                           new_pc_value_mem_stage(19), d(18) => 
                           new_pc_value_mem_stage(18), d(17) => 
                           new_pc_value_mem_stage(17), d(16) => 
                           new_pc_value_mem_stage(16), d(15) => 
                           new_pc_value_mem_stage(15), d(14) => 
                           new_pc_value_mem_stage(14), d(13) => 
                           new_pc_value_mem_stage(13), d(12) => 
                           new_pc_value_mem_stage(12), d(11) => 
                           new_pc_value_mem_stage(11), d(10) => 
                           new_pc_value_mem_stage(10), d(9) => 
                           new_pc_value_mem_stage(9), d(8) => 
                           new_pc_value_mem_stage(8), d(7) => 
                           new_pc_value_mem_stage(7), d(6) => 
                           new_pc_value_mem_stage(6), d(5) => 
                           new_pc_value_mem_stage(5), d(4) => 
                           new_pc_value_mem_stage(4), d(3) => 
                           new_pc_value_mem_stage(3), d(2) => 
                           new_pc_value_mem_stage(2), d(1) => 
                           new_pc_value_mem_stage(1), d(0) => 
                           new_pc_value_mem_stage(0), Q(31) => 
                           IRAM_ADDRESS_31_port, Q(30) => IRAM_ADDRESS_30_port,
                           Q(29) => IRAM_ADDRESS_29_port, Q(28) => 
                           IRAM_ADDRESS_28_port, Q(27) => IRAM_ADDRESS_27_port,
                           Q(26) => IRAM_ADDRESS_26_port, Q(25) => 
                           IRAM_ADDRESS_25_port, Q(24) => IRAM_ADDRESS_24_port,
                           Q(23) => IRAM_ADDRESS_23_port, Q(22) => 
                           IRAM_ADDRESS_22_port, Q(21) => IRAM_ADDRESS_21_port,
                           Q(20) => IRAM_ADDRESS_20_port, Q(19) => 
                           IRAM_ADDRESS_19_port, Q(18) => IRAM_ADDRESS_18_port,
                           Q(17) => IRAM_ADDRESS_17_port, Q(16) => 
                           IRAM_ADDRESS_16_port, Q(15) => IRAM_ADDRESS_15_port,
                           Q(14) => IRAM_ADDRESS_14_port, Q(13) => 
                           IRAM_ADDRESS_13_port, Q(12) => IRAM_ADDRESS_12_port,
                           Q(11) => IRAM_ADDRESS_11_port, Q(10) => 
                           IRAM_ADDRESS_10_port, Q(9) => IRAM_ADDRESS_9_port, 
                           Q(8) => IRAM_ADDRESS_8_port, Q(7) => 
                           IRAM_ADDRESS_7_port, Q(6) => IRAM_ADDRESS_6_port, 
                           Q(5) => IRAM_ADDRESS_5_port, Q(4) => 
                           IRAM_ADDRESS_4_port, Q(3) => IRAM_ADDRESS_3_port, 
                           Q(2) => IRAM_ADDRESS_2_port, Q(1) => 
                           IRAM_ADDRESS_1_port, Q(0) => IRAM_ADDRESS_0_port);
   new_program_counter : reg_nbit_n32_15 port map( clk => clk, reset => 
                           n70_port, d(31) => n2, d(30) => n3, d(29) => n4, 
                           d(28) => n9_port, d(27) => n10_port, d(26) => 
                           n11_port, d(25) => n12_port, d(24) => n13_port, 
                           d(23) => n14_port, d(22) => n15_port, d(21) => 
                           n16_port, d(20) => n17_port, d(19) => n18_port, 
                           d(18) => n19_port, d(17) => n20_port, d(16) => 
                           n21_port, d(15) => n22_port, d(14) => n23_port, 
                           d(13) => n24_port, d(12) => n25_port, d(11) => 
                           n26_port, d(10) => n27_port, d(9) => n28_port, d(8) 
                           => n29_port, d(7) => n30_port, d(6) => n31_port, 
                           d(5) => n32_port, d(4) => n33_port, d(3) => n34_port
                           , d(2) => n35_port, d(1) => n36_port, d(0) => n37, 
                           Q(31) => new_pc_value(31), Q(30) => new_pc_value(30)
                           , Q(29) => new_pc_value(29), Q(28) => 
                           new_pc_value(28), Q(27) => new_pc_value(27), Q(26) 
                           => new_pc_value(26), Q(25) => new_pc_value(25), 
                           Q(24) => new_pc_value(24), Q(23) => new_pc_value(23)
                           , Q(22) => new_pc_value(22), Q(21) => 
                           new_pc_value(21), Q(20) => new_pc_value(20), Q(19) 
                           => new_pc_value(19), Q(18) => new_pc_value(18), 
                           Q(17) => new_pc_value(17), Q(16) => new_pc_value(16)
                           , Q(15) => new_pc_value(15), Q(14) => 
                           new_pc_value(14), Q(13) => new_pc_value(13), Q(12) 
                           => new_pc_value(12), Q(11) => new_pc_value(11), 
                           Q(10) => new_pc_value(10), Q(9) => new_pc_value(9), 
                           Q(8) => new_pc_value(8), Q(7) => new_pc_value(7), 
                           Q(6) => new_pc_value(6), Q(5) => new_pc_value(5), 
                           Q(4) => new_pc_value(4), Q(3) => new_pc_value(3), 
                           Q(2) => new_pc_value(2), Q(1) => new_pc_value(1), 
                           Q(0) => new_pc_value(0));
   instruction_reg : reg_nbit_n32_14 port map( clk => clk, reset => n70_port, 
                           d(31) => n69_port, d(30) => n68_port, d(29) => 
                           n67_port, d(28) => n66_port, d(27) => n65_port, 
                           d(26) => n64_port, d(25) => n63_port, d(24) => 
                           n62_port, d(23) => n61_port, d(22) => n60_port, 
                           d(21) => n59_port, d(20) => n58_port, d(19) => 
                           n57_port, d(18) => n56_port, d(17) => n55_port, 
                           d(16) => n54_port, d(15) => n53_port, d(14) => 
                           n52_port, d(13) => n51_port, d(12) => n50_port, 
                           d(11) => n49_port, d(10) => n48_port, d(9) => 
                           n47_port, d(8) => n46_port, d(7) => n45_port, d(6) 
                           => n44_port, d(5) => n43_port, d(4) => n42_port, 
                           d(3) => n41_port, d(2) => n40_port, d(1) => n39_port
                           , d(0) => n38, Q(31) => curr_instruction_31_port, 
                           Q(30) => curr_instruction_30_port, Q(29) => 
                           curr_instruction_29_port, Q(28) => 
                           curr_instruction_28_port, Q(27) => 
                           curr_instruction_27_port, Q(26) => 
                           curr_instruction_26_port, Q(25) => 
                           curr_instruction_25_port, Q(24) => 
                           curr_instruction_24_port, Q(23) => 
                           curr_instruction_23_port, Q(22) => 
                           curr_instruction_22_port, Q(21) => 
                           curr_instruction_21_port, Q(20) => 
                           curr_instruction_20_port, Q(19) => 
                           curr_instruction_19_port, Q(18) => 
                           curr_instruction_18_port, Q(17) => 
                           curr_instruction_17_port, Q(16) => 
                           curr_instruction_16_port, Q(15) => 
                           curr_instruction_15_port, Q(14) => 
                           curr_instruction_14_port, Q(13) => 
                           curr_instruction_13_port, Q(12) => 
                           curr_instruction_12_port, Q(11) => 
                           curr_instruction_11_port, Q(10) => 
                           curr_instruction_10_port, Q(9) => 
                           curr_instruction_9_port, Q(8) => 
                           curr_instruction_8_port, Q(7) => 
                           curr_instruction_7_port, Q(6) => 
                           curr_instruction_6_port, Q(5) => 
                           curr_instruction_5_port, Q(4) => 
                           curr_instruction_4_port, Q(3) => 
                           curr_instruction_3_port, Q(2) => 
                           curr_instruction_2_port, Q(1) => 
                           curr_instruction_1_port, Q(0) => 
                           curr_instruction_0_port);
   add_79_3_aco : fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_0 port map( A(31) =>
                           IRAM_ADDRESS_31_port, A(30) => IRAM_ADDRESS_30_port,
                           A(29) => IRAM_ADDRESS_29_port, A(28) => 
                           IRAM_ADDRESS_28_port, A(27) => IRAM_ADDRESS_27_port,
                           A(26) => IRAM_ADDRESS_26_port, A(25) => 
                           IRAM_ADDRESS_25_port, A(24) => IRAM_ADDRESS_24_port,
                           A(23) => IRAM_ADDRESS_23_port, A(22) => 
                           IRAM_ADDRESS_22_port, A(21) => IRAM_ADDRESS_21_port,
                           A(20) => IRAM_ADDRESS_20_port, A(19) => 
                           IRAM_ADDRESS_19_port, A(18) => IRAM_ADDRESS_18_port,
                           A(17) => IRAM_ADDRESS_17_port, A(16) => 
                           IRAM_ADDRESS_16_port, A(15) => IRAM_ADDRESS_15_port,
                           A(14) => IRAM_ADDRESS_14_port, A(13) => 
                           IRAM_ADDRESS_13_port, A(12) => IRAM_ADDRESS_12_port,
                           A(11) => IRAM_ADDRESS_11_port, A(10) => 
                           IRAM_ADDRESS_10_port, A(9) => IRAM_ADDRESS_9_port, 
                           A(8) => IRAM_ADDRESS_8_port, A(7) => 
                           IRAM_ADDRESS_7_port, A(6) => IRAM_ADDRESS_6_port, 
                           A(5) => IRAM_ADDRESS_5_port, A(4) => 
                           IRAM_ADDRESS_4_port, A(3) => IRAM_ADDRESS_3_port, 
                           A(2) => IRAM_ADDRESS_2_port, A(1) => 
                           IRAM_ADDRESS_1_port, A(0) => IRAM_ADDRESS_0_port, 
                           B(31) => n7_port, B(30) => n7_port, B(29) => n7_port
                           , B(28) => n7_port, B(27) => n7_port, B(26) => 
                           n7_port, B(25) => n7_port, B(24) => n7_port, B(23) 
                           => n7_port, B(22) => n7_port, B(21) => n7_port, 
                           B(20) => n7_port, B(19) => n7_port, B(18) => n7_port
                           , B(17) => n7_port, B(16) => n7_port, B(15) => 
                           n7_port, B(14) => n7_port, B(13) => n7_port, B(12) 
                           => n7_port, B(11) => n7_port, B(10) => n7_port, B(9)
                           => n7_port, B(8) => n7_port, B(7) => n7_port, B(6) 
                           => n7_port, B(5) => n7_port, B(4) => n7_port, B(3) 
                           => n7_port, B(2) => iram_enable_cu, B(1) => n5_port,
                           B(0) => n5_port, CI => n7_port, SUM(31) => N70, 
                           SUM(30) => N69, SUM(29) => N68, SUM(28) => N67, 
                           SUM(27) => N66, SUM(26) => N65, SUM(25) => N64, 
                           SUM(24) => N63, SUM(23) => N62, SUM(22) => N61, 
                           SUM(21) => N60, SUM(20) => N59, SUM(19) => N58, 
                           SUM(18) => N57, SUM(17) => N56, SUM(16) => N55, 
                           SUM(15) => N54, SUM(14) => N53, SUM(13) => N52, 
                           SUM(12) => N51, SUM(11) => N50, SUM(10) => N49, 
                           SUM(9) => N48, SUM(8) => N47, SUM(7) => N46, SUM(6) 
                           => N45, SUM(5) => N44, SUM(4) => N43, SUM(3) => N42,
                           SUM(2) => N41, SUM(1) => N40, SUM(0) => N39, CO => 
                           n_5534);
   add_79 : fetch_stage_IR_SIZE32_PC_SIZE32_DW01_add_1 port map( A(31) => 
                           new_pc_value_mem_stage(31), A(30) => 
                           new_pc_value_mem_stage(30), A(29) => 
                           new_pc_value_mem_stage(29), A(28) => 
                           new_pc_value_mem_stage(28), A(27) => 
                           new_pc_value_mem_stage(27), A(26) => 
                           new_pc_value_mem_stage(26), A(25) => 
                           new_pc_value_mem_stage(25), A(24) => 
                           new_pc_value_mem_stage(24), A(23) => 
                           new_pc_value_mem_stage(23), A(22) => 
                           new_pc_value_mem_stage(22), A(21) => 
                           new_pc_value_mem_stage(21), A(20) => 
                           new_pc_value_mem_stage(20), A(19) => 
                           new_pc_value_mem_stage(19), A(18) => 
                           new_pc_value_mem_stage(18), A(17) => 
                           new_pc_value_mem_stage(17), A(16) => 
                           new_pc_value_mem_stage(16), A(15) => 
                           new_pc_value_mem_stage(15), A(14) => 
                           new_pc_value_mem_stage(14), A(13) => 
                           new_pc_value_mem_stage(13), A(12) => 
                           new_pc_value_mem_stage(12), A(11) => 
                           new_pc_value_mem_stage(11), A(10) => 
                           new_pc_value_mem_stage(10), A(9) => 
                           new_pc_value_mem_stage(9), A(8) => 
                           new_pc_value_mem_stage(8), A(7) => 
                           new_pc_value_mem_stage(7), A(6) => 
                           new_pc_value_mem_stage(6), A(5) => 
                           new_pc_value_mem_stage(5), A(4) => 
                           new_pc_value_mem_stage(4), A(3) => 
                           new_pc_value_mem_stage(3), A(2) => 
                           new_pc_value_mem_stage(2), A(1) => 
                           new_pc_value_mem_stage(1), A(0) => 
                           new_pc_value_mem_stage(0), B(31) => n8_port, B(30) 
                           => n8_port, B(29) => n8_port, B(28) => n8_port, 
                           B(27) => n8_port, B(26) => n8_port, B(25) => n8_port
                           , B(24) => n8_port, B(23) => n8_port, B(22) => 
                           n8_port, B(21) => n8_port, B(20) => n8_port, B(19) 
                           => n8_port, B(18) => n8_port, B(17) => n8_port, 
                           B(16) => n8_port, B(15) => n8_port, B(14) => n8_port
                           , B(13) => n8_port, B(12) => n8_port, B(11) => 
                           n8_port, B(10) => n8_port, B(9) => n8_port, B(8) => 
                           n8_port, B(7) => n8_port, B(6) => n8_port, B(5) => 
                           n8_port, B(4) => n8_port, B(3) => n8_port, B(2) => 
                           n6_port, B(1) => n5_port, B(0) => n5_port, CI => 
                           n8_port, SUM(31) => N36, SUM(30) => N35, SUM(29) => 
                           N34, SUM(28) => N33, SUM(27) => N32, SUM(26) => N31,
                           SUM(25) => N30, SUM(24) => N29, SUM(23) => N28, 
                           SUM(22) => N27, SUM(21) => N26, SUM(20) => N25, 
                           SUM(19) => N24, SUM(18) => N23, SUM(17) => N22, 
                           SUM(16) => N21, SUM(15) => N20, SUM(14) => N19, 
                           SUM(13) => N18, SUM(12) => N17, SUM(11) => N16, 
                           SUM(10) => N15, SUM(9) => N14, SUM(8) => N13, SUM(7)
                           => N12, SUM(6) => N11, SUM(5) => N10, SUM(4) => N9, 
                           SUM(3) => N8, SUM(2) => N7, SUM(1) => N6, SUM(0) => 
                           N5, CO => n_5535);
   U5 : INV_X8 port map( A => rst, ZN => n70_port);
   U6 : NOR2_X4 port map( A1 => update_pc_branch, A2 => branch_taken, ZN => n1)
                           ;
   U9 : MUX2_X1 port map( A => N36, B => N70, S => n1, Z => n2);
   U10 : MUX2_X1 port map( A => N35, B => N69, S => n1, Z => n3);
   U11 : MUX2_X1 port map( A => N34, B => N68, S => n1, Z => n4);
   U12 : MUX2_X1 port map( A => N33, B => N67, S => n1, Z => n9_port);
   U13 : MUX2_X1 port map( A => N32, B => N66, S => n1, Z => n10_port);
   U14 : MUX2_X1 port map( A => N31, B => N65, S => n1, Z => n11_port);
   U15 : MUX2_X1 port map( A => N30, B => N64, S => n1, Z => n12_port);
   U16 : MUX2_X1 port map( A => N29, B => N63, S => n1, Z => n13_port);
   U17 : MUX2_X1 port map( A => N28, B => N62, S => n1, Z => n14_port);
   U18 : MUX2_X1 port map( A => N27, B => N61, S => n1, Z => n15_port);
   U19 : MUX2_X1 port map( A => N26, B => N60, S => n1, Z => n16_port);
   U20 : MUX2_X1 port map( A => N25, B => N59, S => n1, Z => n17_port);
   U21 : MUX2_X1 port map( A => N24, B => N58, S => n1, Z => n18_port);
   U22 : MUX2_X1 port map( A => N23, B => N57, S => n1, Z => n19_port);
   U23 : MUX2_X1 port map( A => N22, B => N56, S => n1, Z => n20_port);
   U24 : MUX2_X1 port map( A => N21, B => N55, S => n1, Z => n21_port);
   U25 : MUX2_X1 port map( A => N20, B => N54, S => n1, Z => n22_port);
   U26 : MUX2_X1 port map( A => N19, B => N53, S => n1, Z => n23_port);
   U27 : MUX2_X1 port map( A => N18, B => N52, S => n1, Z => n24_port);
   U28 : MUX2_X1 port map( A => N17, B => N51, S => n1, Z => n25_port);
   U29 : MUX2_X1 port map( A => N16, B => N50, S => n1, Z => n26_port);
   U30 : MUX2_X1 port map( A => N15, B => N49, S => n1, Z => n27_port);
   U31 : MUX2_X1 port map( A => N14, B => N48, S => n1, Z => n28_port);
   U32 : MUX2_X1 port map( A => N13, B => N47, S => n1, Z => n29_port);
   U33 : MUX2_X1 port map( A => N12, B => N46, S => n1, Z => n30_port);
   U34 : MUX2_X1 port map( A => N11, B => N45, S => n1, Z => n31_port);
   U35 : MUX2_X1 port map( A => N10, B => N44, S => n1, Z => n32_port);
   U36 : MUX2_X1 port map( A => N9, B => N43, S => n1, Z => n33_port);
   U37 : MUX2_X1 port map( A => N8, B => N42, S => n1, Z => n34_port);
   U38 : MUX2_X1 port map( A => N7, B => N41, S => n1, Z => n35_port);
   U39 : MUX2_X1 port map( A => N6, B => N40, S => n1, Z => n36_port);
   U40 : MUX2_X1 port map( A => N5, B => N39, S => n1, Z => n37);
   U41 : MUX2_X1 port map( A => IRAM_DATA(31), B => curr_instruction_0_port, S 
                           => stall, Z => n38);
   U42 : MUX2_X1 port map( A => IRAM_DATA(30), B => curr_instruction_1_port, S 
                           => stall, Z => n39_port);
   U43 : MUX2_X1 port map( A => IRAM_DATA(29), B => curr_instruction_2_port, S 
                           => stall, Z => n40_port);
   U44 : MUX2_X1 port map( A => IRAM_DATA(28), B => curr_instruction_3_port, S 
                           => stall, Z => n41_port);
   U45 : MUX2_X1 port map( A => IRAM_DATA(27), B => curr_instruction_4_port, S 
                           => stall, Z => n42_port);
   U46 : MUX2_X1 port map( A => IRAM_DATA(26), B => curr_instruction_5_port, S 
                           => stall, Z => n43_port);
   U47 : MUX2_X1 port map( A => IRAM_DATA(25), B => curr_instruction_6_port, S 
                           => stall, Z => n44_port);
   U48 : MUX2_X1 port map( A => IRAM_DATA(24), B => curr_instruction_7_port, S 
                           => stall, Z => n45_port);
   U49 : MUX2_X1 port map( A => IRAM_DATA(23), B => curr_instruction_8_port, S 
                           => stall, Z => n46_port);
   U50 : MUX2_X1 port map( A => IRAM_DATA(22), B => curr_instruction_9_port, S 
                           => stall, Z => n47_port);
   U51 : MUX2_X1 port map( A => IRAM_DATA(21), B => curr_instruction_10_port, S
                           => stall, Z => n48_port);
   U52 : MUX2_X1 port map( A => IRAM_DATA(20), B => curr_instruction_11_port, S
                           => stall, Z => n49_port);
   U53 : MUX2_X1 port map( A => IRAM_DATA(19), B => curr_instruction_12_port, S
                           => stall, Z => n50_port);
   U54 : MUX2_X1 port map( A => IRAM_DATA(18), B => curr_instruction_13_port, S
                           => stall, Z => n51_port);
   U55 : MUX2_X1 port map( A => IRAM_DATA(17), B => curr_instruction_14_port, S
                           => stall, Z => n52_port);
   U56 : MUX2_X1 port map( A => IRAM_DATA(16), B => curr_instruction_15_port, S
                           => stall, Z => n53_port);
   U57 : MUX2_X1 port map( A => IRAM_DATA(15), B => curr_instruction_16_port, S
                           => stall, Z => n54_port);
   U58 : MUX2_X1 port map( A => IRAM_DATA(14), B => curr_instruction_17_port, S
                           => stall, Z => n55_port);
   U59 : MUX2_X1 port map( A => IRAM_DATA(13), B => curr_instruction_18_port, S
                           => stall, Z => n56_port);
   U60 : MUX2_X1 port map( A => IRAM_DATA(12), B => curr_instruction_19_port, S
                           => stall, Z => n57_port);
   U61 : MUX2_X1 port map( A => IRAM_DATA(11), B => curr_instruction_20_port, S
                           => stall, Z => n58_port);
   U62 : MUX2_X1 port map( A => IRAM_DATA(10), B => curr_instruction_21_port, S
                           => stall, Z => n59_port);
   U63 : MUX2_X1 port map( A => IRAM_DATA(9), B => curr_instruction_22_port, S 
                           => stall, Z => n60_port);
   U64 : MUX2_X1 port map( A => IRAM_DATA(8), B => curr_instruction_23_port, S 
                           => stall, Z => n61_port);
   U65 : MUX2_X1 port map( A => IRAM_DATA(7), B => curr_instruction_24_port, S 
                           => stall, Z => n62_port);
   U66 : MUX2_X1 port map( A => IRAM_DATA(6), B => curr_instruction_25_port, S 
                           => stall, Z => n63_port);
   U67 : MUX2_X1 port map( A => IRAM_DATA(5), B => curr_instruction_26_port, S 
                           => stall, Z => n64_port);
   U68 : MUX2_X1 port map( A => IRAM_DATA(4), B => curr_instruction_27_port, S 
                           => stall, Z => n65_port);
   U69 : MUX2_X1 port map( A => IRAM_DATA(3), B => curr_instruction_28_port, S 
                           => stall, Z => n66_port);
   U70 : MUX2_X1 port map( A => IRAM_DATA(2), B => curr_instruction_29_port, S 
                           => stall, Z => n67_port);
   U71 : MUX2_X1 port map( A => IRAM_DATA(1), B => curr_instruction_30_port, S 
                           => stall, Z => n68_port);
   U72 : MUX2_X1 port map( A => IRAM_DATA(0), B => curr_instruction_31_port, S 
                           => stall, Z => n69_port);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity reg_nbit_n22_0 is

   port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0);  Q 
         : out std_logic_vector (21 downto 0));

end reg_nbit_n22_0;

architecture SYN_struc of reg_nbit_n22_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FD_2229
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2230
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2231
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2232
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2233
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2234
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2235
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2236
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2237
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2238
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2239
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2240
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2241
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2242
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2243
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2244
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2245
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2246
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2247
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2248
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2249
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_0
      port( D, CK, RESET : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   D_I_0 : FD_0 port map( D => d(0), CK => n1, RESET => reset, Q => Q(0));
   D_I_1 : FD_2249 port map( D => d(1), CK => n2, RESET => reset, Q => Q(1));
   D_I_2 : FD_2248 port map( D => d(2), CK => n2, RESET => reset, Q => Q(2));
   D_I_3 : FD_2247 port map( D => d(3), CK => n2, RESET => reset, Q => Q(3));
   D_I_4 : FD_2246 port map( D => d(4), CK => n2, RESET => reset, Q => Q(4));
   D_I_5 : FD_2245 port map( D => d(5), CK => n2, RESET => reset, Q => Q(5));
   D_I_6 : FD_2244 port map( D => d(6), CK => n2, RESET => reset, Q => Q(6));
   D_I_7 : FD_2243 port map( D => d(7), CK => n2, RESET => reset, Q => Q(7));
   D_I_8 : FD_2242 port map( D => d(8), CK => n2, RESET => reset, Q => Q(8));
   D_I_9 : FD_2241 port map( D => d(9), CK => n2, RESET => reset, Q => Q(9));
   D_I_10 : FD_2240 port map( D => d(10), CK => n2, RESET => reset, Q => Q(10))
                           ;
   D_I_11 : FD_2239 port map( D => d(11), CK => n2, RESET => reset, Q => Q(11))
                           ;
   D_I_12 : FD_2238 port map( D => d(12), CK => n1, RESET => reset, Q => Q(12))
                           ;
   D_I_13 : FD_2237 port map( D => d(13), CK => n1, RESET => reset, Q => Q(13))
                           ;
   D_I_14 : FD_2236 port map( D => d(14), CK => n1, RESET => reset, Q => Q(14))
                           ;
   D_I_15 : FD_2235 port map( D => d(15), CK => n1, RESET => reset, Q => Q(15))
                           ;
   D_I_16 : FD_2234 port map( D => d(16), CK => n1, RESET => reset, Q => Q(16))
                           ;
   D_I_17 : FD_2233 port map( D => d(17), CK => n1, RESET => reset, Q => Q(17))
                           ;
   D_I_18 : FD_2232 port map( D => d(18), CK => n1, RESET => reset, Q => Q(18))
                           ;
   D_I_19 : FD_2231 port map( D => d(19), CK => n1, RESET => reset, Q => Q(19))
                           ;
   D_I_20 : FD_2230 port map( D => d(20), CK => n1, RESET => reset, Q => Q(20))
                           ;
   D_I_21 : FD_2229 port map( D => d(21), CK => n1, RESET => reset, Q => Q(21))
                           ;
   U1 : BUF_X1 port map( A => clk, Z => n2);
   U2 : BUF_X1 port map( A => clk, Z => n1);

end SYN_struc;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPATH_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 is

   port( clk, rst : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0);  iram_enable_cu : in std_logic;  
         iram_ready_cu : out std_logic;  stall : in std_logic;  
         curr_instruction_to_cu : out std_logic_vector (31 downto 0);  
         enable_rf, read_rf_p1, read_rf_p2, write_rf, rtype_itypen, 
         compute_sext, jump_sext : in std_logic;  alu_op_type : in 
         std_logic_vector (3 downto 0);  sel_val_a, sel_val_b, signed_notsigned
         : in std_logic;  evaluate_branch : in std_logic_vector (1 downto 0);  
         alu_cin : in std_logic;  alu_overflow, zero_mul_detect, mul_exeception
         : out std_logic;  dram_enable_cu, dram_r_nw_cu : in std_logic;  
         dram_ready_cu : out std_logic;  update_pc_branch, select_wb : in 
         std_logic);

end DATAPATH_N32_RF_REGS32_IR_SIZE32_PC_SIZE32;

architecture SYN_structural of DATAPATH_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 is

   component write_back_stage_N32
      port( data_from_memory, data_from_alu : in std_logic_vector (31 downto 0)
            ;  data_to_rf : out std_logic_vector (31 downto 0);  select_wb : in
            std_logic);
   end component;
   
   component memory_stage_N32_PC_SIZE32
      port( clk, rst : in std_logic;  new_pc_value : in std_logic_vector (31 
            downto 0);  new_pc_value_branch : out std_logic_vector (31 downto 
            0);  select_pc : in std_logic;  alu_output_val, value_to_mem : in 
            std_logic_vector (31 downto 0);  data_from_memory, data_from_alu : 
            out std_logic_vector (31 downto 0);  dram_enable_cu, dram_r_nw_cu :
            in std_logic;  dram_ready_cu : out std_logic;  DRAM_ADDRESS : out 
            std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : 
            out std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
            std_logic_vector (31 downto 0));
   end component;
   
   component execute_stage_N32_PC_SIZE32
      port( clk, rst : in std_logic;  val_a, val_b, val_immediate, 
            new_prog_counter_val_exe : in std_logic_vector (31 downto 0);  
            branch_condition : out std_logic;  prog_counter_forwaded, 
            alu_output_val, value_to_mem : out std_logic_vector (31 downto 0); 
            signed_notsigned : in std_logic;  alu_op_type : in std_logic_vector
            (3 downto 0);  sel_val_a, sel_val_b, cin : in std_logic;  overflow,
            zero_mul_detect, mul_exeception : out std_logic;  evaluate_branch :
            in std_logic_vector (1 downto 0));
   end component;
   
   component decode_stage_N32_RF_REGS32_IR_SIZE32_PC_SIZE32
      port( clk, rst : in std_logic;  new_prog_counter_val, instruction_reg : 
            in std_logic_vector (31 downto 0);  val_a, new_prog_counter_val_exe
            , val_b, val_immediate : out std_logic_vector (31 downto 0);  
            update_reg_value : in std_logic_vector (31 downto 0);  enable_rf, 
            read_rf_p1, read_rf_p2, write_rf, rtype_itypen, jump_sext, 
            compute_sext : in std_logic);
   end component;
   
   component fetch_stage_IR_SIZE32_PC_SIZE32
      port( clk, rst : in std_logic;  new_pc_value_mem_stage : in 
            std_logic_vector (31 downto 0);  branch_taken : in std_logic;  
            new_pc_value, IRAM_ADDRESS : out std_logic_vector (31 downto 0);  
            IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  IRAM_DATA
            : in std_logic_vector (0 to 31);  curr_instruction : out 
            std_logic_vector (31 downto 0);  iram_enable_cu, update_pc_branch, 
            stall : in std_logic;  iram_ready_cu : out std_logic);
   end component;
   
   signal curr_instruction_to_cu_31_port, curr_instruction_to_cu_30_port, 
      curr_instruction_to_cu_29_port, curr_instruction_to_cu_28_port, 
      curr_instruction_to_cu_27_port, curr_instruction_to_cu_26_port, 
      curr_instruction_to_cu_25_port, curr_instruction_to_cu_24_port, 
      curr_instruction_to_cu_23_port, curr_instruction_to_cu_22_port, 
      curr_instruction_to_cu_21_port, curr_instruction_to_cu_20_port, 
      curr_instruction_to_cu_19_port, curr_instruction_to_cu_18_port, 
      curr_instruction_to_cu_17_port, curr_instruction_to_cu_16_port, 
      curr_instruction_to_cu_15_port, curr_instruction_to_cu_14_port, 
      curr_instruction_to_cu_13_port, curr_instruction_to_cu_12_port, 
      curr_instruction_to_cu_11_port, curr_instruction_to_cu_10_port, 
      curr_instruction_to_cu_9_port, curr_instruction_to_cu_8_port, 
      curr_instruction_to_cu_7_port, curr_instruction_to_cu_6_port, 
      curr_instruction_to_cu_5_port, curr_instruction_to_cu_4_port, 
      curr_instruction_to_cu_3_port, curr_instruction_to_cu_2_port, 
      curr_instruction_to_cu_1_port, curr_instruction_to_cu_0_port, 
      new_pc_value_mem_stage_i_31_port, new_pc_value_mem_stage_i_30_port, 
      new_pc_value_mem_stage_i_29_port, new_pc_value_mem_stage_i_28_port, 
      new_pc_value_mem_stage_i_27_port, new_pc_value_mem_stage_i_26_port, 
      new_pc_value_mem_stage_i_25_port, new_pc_value_mem_stage_i_24_port, 
      new_pc_value_mem_stage_i_23_port, new_pc_value_mem_stage_i_22_port, 
      new_pc_value_mem_stage_i_21_port, new_pc_value_mem_stage_i_20_port, 
      new_pc_value_mem_stage_i_19_port, new_pc_value_mem_stage_i_18_port, 
      new_pc_value_mem_stage_i_17_port, new_pc_value_mem_stage_i_16_port, 
      new_pc_value_mem_stage_i_15_port, new_pc_value_mem_stage_i_14_port, 
      new_pc_value_mem_stage_i_13_port, new_pc_value_mem_stage_i_12_port, 
      new_pc_value_mem_stage_i_11_port, new_pc_value_mem_stage_i_10_port, 
      new_pc_value_mem_stage_i_9_port, new_pc_value_mem_stage_i_8_port, 
      new_pc_value_mem_stage_i_7_port, new_pc_value_mem_stage_i_6_port, 
      new_pc_value_mem_stage_i_5_port, new_pc_value_mem_stage_i_4_port, 
      new_pc_value_mem_stage_i_3_port, new_pc_value_mem_stage_i_2_port, 
      new_pc_value_mem_stage_i_1_port, new_pc_value_mem_stage_i_0_port, 
      branch_condition_i_0_port, new_pc_value_decode_31_port, 
      new_pc_value_decode_30_port, new_pc_value_decode_29_port, 
      new_pc_value_decode_28_port, new_pc_value_decode_27_port, 
      new_pc_value_decode_26_port, new_pc_value_decode_25_port, 
      new_pc_value_decode_24_port, new_pc_value_decode_23_port, 
      new_pc_value_decode_22_port, new_pc_value_decode_21_port, 
      new_pc_value_decode_20_port, new_pc_value_decode_19_port, 
      new_pc_value_decode_18_port, new_pc_value_decode_17_port, 
      new_pc_value_decode_16_port, new_pc_value_decode_15_port, 
      new_pc_value_decode_14_port, new_pc_value_decode_13_port, 
      new_pc_value_decode_12_port, new_pc_value_decode_11_port, 
      new_pc_value_decode_10_port, new_pc_value_decode_9_port, 
      new_pc_value_decode_8_port, new_pc_value_decode_7_port, 
      new_pc_value_decode_6_port, new_pc_value_decode_5_port, 
      new_pc_value_decode_4_port, new_pc_value_decode_3_port, 
      new_pc_value_decode_2_port, new_pc_value_decode_1_port, 
      new_pc_value_decode_0_port, val_a_i_31_port, val_a_i_30_port, 
      val_a_i_29_port, val_a_i_28_port, val_a_i_27_port, val_a_i_26_port, 
      val_a_i_25_port, val_a_i_24_port, val_a_i_23_port, val_a_i_22_port, 
      val_a_i_21_port, val_a_i_20_port, val_a_i_19_port, val_a_i_18_port, 
      val_a_i_17_port, val_a_i_16_port, val_a_i_15_port, val_a_i_14_port, 
      val_a_i_13_port, val_a_i_12_port, val_a_i_11_port, val_a_i_10_port, 
      val_a_i_9_port, val_a_i_8_port, val_a_i_7_port, val_a_i_6_port, 
      val_a_i_5_port, val_a_i_4_port, val_a_i_3_port, val_a_i_2_port, 
      val_a_i_1_port, val_a_i_0_port, new_prog_counter_val_exe_i_31_port, 
      new_prog_counter_val_exe_i_30_port, new_prog_counter_val_exe_i_29_port, 
      new_prog_counter_val_exe_i_28_port, new_prog_counter_val_exe_i_27_port, 
      new_prog_counter_val_exe_i_26_port, new_prog_counter_val_exe_i_25_port, 
      new_prog_counter_val_exe_i_24_port, new_prog_counter_val_exe_i_23_port, 
      new_prog_counter_val_exe_i_22_port, new_prog_counter_val_exe_i_21_port, 
      new_prog_counter_val_exe_i_20_port, new_prog_counter_val_exe_i_19_port, 
      new_prog_counter_val_exe_i_18_port, new_prog_counter_val_exe_i_17_port, 
      new_prog_counter_val_exe_i_16_port, new_prog_counter_val_exe_i_15_port, 
      new_prog_counter_val_exe_i_14_port, new_prog_counter_val_exe_i_13_port, 
      new_prog_counter_val_exe_i_12_port, new_prog_counter_val_exe_i_11_port, 
      new_prog_counter_val_exe_i_10_port, new_prog_counter_val_exe_i_9_port, 
      new_prog_counter_val_exe_i_8_port, new_prog_counter_val_exe_i_7_port, 
      new_prog_counter_val_exe_i_6_port, new_prog_counter_val_exe_i_5_port, 
      new_prog_counter_val_exe_i_4_port, new_prog_counter_val_exe_i_3_port, 
      new_prog_counter_val_exe_i_2_port, new_prog_counter_val_exe_i_1_port, 
      new_prog_counter_val_exe_i_0_port, val_b_i_31_port, val_b_i_30_port, 
      val_b_i_29_port, val_b_i_28_port, val_b_i_27_port, val_b_i_26_port, 
      val_b_i_25_port, val_b_i_24_port, val_b_i_23_port, val_b_i_22_port, 
      val_b_i_21_port, val_b_i_20_port, val_b_i_19_port, val_b_i_18_port, 
      val_b_i_17_port, val_b_i_16_port, val_b_i_15_port, val_b_i_14_port, 
      val_b_i_13_port, val_b_i_12_port, val_b_i_11_port, val_b_i_10_port, 
      val_b_i_9_port, val_b_i_8_port, val_b_i_7_port, val_b_i_6_port, 
      val_b_i_5_port, val_b_i_4_port, val_b_i_3_port, val_b_i_2_port, 
      val_b_i_1_port, val_b_i_0_port, val_immediate_i_31_port, 
      val_immediate_i_30_port, val_immediate_i_29_port, val_immediate_i_28_port
      , val_immediate_i_27_port, val_immediate_i_26_port, 
      val_immediate_i_25_port, val_immediate_i_24_port, val_immediate_i_23_port
      , val_immediate_i_22_port, val_immediate_i_21_port, 
      val_immediate_i_20_port, val_immediate_i_19_port, val_immediate_i_18_port
      , val_immediate_i_17_port, val_immediate_i_16_port, 
      val_immediate_i_15_port, val_immediate_i_14_port, val_immediate_i_13_port
      , val_immediate_i_12_port, val_immediate_i_11_port, 
      val_immediate_i_10_port, val_immediate_i_9_port, val_immediate_i_8_port, 
      val_immediate_i_7_port, val_immediate_i_6_port, val_immediate_i_5_port, 
      val_immediate_i_4_port, val_immediate_i_3_port, val_immediate_i_2_port, 
      val_immediate_i_1_port, val_immediate_i_0_port, 
      update_reg_value_i_31_port, update_reg_value_i_30_port, 
      update_reg_value_i_29_port, update_reg_value_i_28_port, 
      update_reg_value_i_27_port, update_reg_value_i_26_port, 
      update_reg_value_i_25_port, update_reg_value_i_24_port, 
      update_reg_value_i_23_port, update_reg_value_i_22_port, 
      update_reg_value_i_21_port, update_reg_value_i_20_port, 
      update_reg_value_i_19_port, update_reg_value_i_18_port, 
      update_reg_value_i_17_port, update_reg_value_i_16_port, 
      update_reg_value_i_15_port, update_reg_value_i_14_port, 
      update_reg_value_i_13_port, update_reg_value_i_12_port, 
      update_reg_value_i_11_port, update_reg_value_i_10_port, 
      update_reg_value_i_9_port, update_reg_value_i_8_port, 
      update_reg_value_i_7_port, update_reg_value_i_6_port, 
      update_reg_value_i_5_port, update_reg_value_i_4_port, 
      update_reg_value_i_3_port, update_reg_value_i_2_port, 
      update_reg_value_i_1_port, update_reg_value_i_0_port, 
      prog_counter_forwaded_i_31_port, prog_counter_forwaded_i_30_port, 
      prog_counter_forwaded_i_29_port, prog_counter_forwaded_i_28_port, 
      prog_counter_forwaded_i_27_port, prog_counter_forwaded_i_26_port, 
      prog_counter_forwaded_i_25_port, prog_counter_forwaded_i_24_port, 
      prog_counter_forwaded_i_23_port, prog_counter_forwaded_i_22_port, 
      prog_counter_forwaded_i_21_port, prog_counter_forwaded_i_20_port, 
      prog_counter_forwaded_i_19_port, prog_counter_forwaded_i_18_port, 
      prog_counter_forwaded_i_17_port, prog_counter_forwaded_i_16_port, 
      prog_counter_forwaded_i_15_port, prog_counter_forwaded_i_14_port, 
      prog_counter_forwaded_i_13_port, prog_counter_forwaded_i_12_port, 
      prog_counter_forwaded_i_11_port, prog_counter_forwaded_i_10_port, 
      prog_counter_forwaded_i_9_port, prog_counter_forwaded_i_8_port, 
      prog_counter_forwaded_i_7_port, prog_counter_forwaded_i_6_port, 
      prog_counter_forwaded_i_5_port, prog_counter_forwaded_i_4_port, 
      prog_counter_forwaded_i_3_port, prog_counter_forwaded_i_2_port, 
      prog_counter_forwaded_i_1_port, prog_counter_forwaded_i_0_port, 
      alu_output_val_i_31_port, alu_output_val_i_30_port, 
      alu_output_val_i_29_port, alu_output_val_i_28_port, 
      alu_output_val_i_27_port, alu_output_val_i_26_port, 
      alu_output_val_i_25_port, alu_output_val_i_24_port, 
      alu_output_val_i_23_port, alu_output_val_i_22_port, 
      alu_output_val_i_21_port, alu_output_val_i_20_port, 
      alu_output_val_i_19_port, alu_output_val_i_18_port, 
      alu_output_val_i_17_port, alu_output_val_i_16_port, 
      alu_output_val_i_15_port, alu_output_val_i_14_port, 
      alu_output_val_i_13_port, alu_output_val_i_12_port, 
      alu_output_val_i_11_port, alu_output_val_i_10_port, 
      alu_output_val_i_9_port, alu_output_val_i_8_port, alu_output_val_i_7_port
      , alu_output_val_i_6_port, alu_output_val_i_5_port, 
      alu_output_val_i_4_port, alu_output_val_i_3_port, alu_output_val_i_2_port
      , alu_output_val_i_1_port, alu_output_val_i_0_port, 
      value_to_mem_i_31_port, value_to_mem_i_30_port, value_to_mem_i_29_port, 
      value_to_mem_i_28_port, value_to_mem_i_27_port, value_to_mem_i_26_port, 
      value_to_mem_i_25_port, value_to_mem_i_24_port, value_to_mem_i_23_port, 
      value_to_mem_i_22_port, value_to_mem_i_21_port, value_to_mem_i_20_port, 
      value_to_mem_i_19_port, value_to_mem_i_18_port, value_to_mem_i_17_port, 
      value_to_mem_i_16_port, value_to_mem_i_15_port, value_to_mem_i_14_port, 
      value_to_mem_i_13_port, value_to_mem_i_12_port, value_to_mem_i_11_port, 
      value_to_mem_i_10_port, value_to_mem_i_9_port, value_to_mem_i_8_port, 
      value_to_mem_i_7_port, value_to_mem_i_6_port, value_to_mem_i_5_port, 
      value_to_mem_i_4_port, value_to_mem_i_3_port, value_to_mem_i_2_port, 
      value_to_mem_i_1_port, value_to_mem_i_0_port, data_from_memory_i_31_port,
      data_from_memory_i_30_port, data_from_memory_i_29_port, 
      data_from_memory_i_28_port, data_from_memory_i_27_port, 
      data_from_memory_i_26_port, data_from_memory_i_25_port, 
      data_from_memory_i_24_port, data_from_memory_i_23_port, 
      data_from_memory_i_22_port, data_from_memory_i_21_port, 
      data_from_memory_i_20_port, data_from_memory_i_19_port, 
      data_from_memory_i_18_port, data_from_memory_i_17_port, 
      data_from_memory_i_16_port, data_from_memory_i_15_port, 
      data_from_memory_i_14_port, data_from_memory_i_13_port, 
      data_from_memory_i_12_port, data_from_memory_i_11_port, 
      data_from_memory_i_10_port, data_from_memory_i_9_port, 
      data_from_memory_i_8_port, data_from_memory_i_7_port, 
      data_from_memory_i_6_port, data_from_memory_i_5_port, 
      data_from_memory_i_4_port, data_from_memory_i_3_port, 
      data_from_memory_i_2_port, data_from_memory_i_1_port, 
      data_from_memory_i_0_port, data_from_alu_i_31_port, 
      data_from_alu_i_30_port, data_from_alu_i_29_port, data_from_alu_i_28_port
      , data_from_alu_i_27_port, data_from_alu_i_26_port, 
      data_from_alu_i_25_port, data_from_alu_i_24_port, data_from_alu_i_23_port
      , data_from_alu_i_22_port, data_from_alu_i_21_port, 
      data_from_alu_i_20_port, data_from_alu_i_19_port, data_from_alu_i_18_port
      , data_from_alu_i_17_port, data_from_alu_i_16_port, 
      data_from_alu_i_15_port, data_from_alu_i_14_port, data_from_alu_i_13_port
      , data_from_alu_i_12_port, data_from_alu_i_11_port, 
      data_from_alu_i_10_port, data_from_alu_i_9_port, data_from_alu_i_8_port, 
      data_from_alu_i_7_port, data_from_alu_i_6_port, data_from_alu_i_5_port, 
      data_from_alu_i_4_port, data_from_alu_i_3_port, data_from_alu_i_2_port, 
      data_from_alu_i_1_port, data_from_alu_i_0_port, n_5536, n_5537 : 
      std_logic;

begin
   curr_instruction_to_cu <= ( curr_instruction_to_cu_31_port, 
      curr_instruction_to_cu_30_port, curr_instruction_to_cu_29_port, 
      curr_instruction_to_cu_28_port, curr_instruction_to_cu_27_port, 
      curr_instruction_to_cu_26_port, curr_instruction_to_cu_25_port, 
      curr_instruction_to_cu_24_port, curr_instruction_to_cu_23_port, 
      curr_instruction_to_cu_22_port, curr_instruction_to_cu_21_port, 
      curr_instruction_to_cu_20_port, curr_instruction_to_cu_19_port, 
      curr_instruction_to_cu_18_port, curr_instruction_to_cu_17_port, 
      curr_instruction_to_cu_16_port, curr_instruction_to_cu_15_port, 
      curr_instruction_to_cu_14_port, curr_instruction_to_cu_13_port, 
      curr_instruction_to_cu_12_port, curr_instruction_to_cu_11_port, 
      curr_instruction_to_cu_10_port, curr_instruction_to_cu_9_port, 
      curr_instruction_to_cu_8_port, curr_instruction_to_cu_7_port, 
      curr_instruction_to_cu_6_port, curr_instruction_to_cu_5_port, 
      curr_instruction_to_cu_4_port, curr_instruction_to_cu_3_port, 
      curr_instruction_to_cu_2_port, curr_instruction_to_cu_1_port, 
      curr_instruction_to_cu_0_port );
   
   fetch_stage_dp : fetch_stage_IR_SIZE32_PC_SIZE32 port map( clk => clk, rst 
                           => rst, new_pc_value_mem_stage(31) => 
                           new_pc_value_mem_stage_i_31_port, 
                           new_pc_value_mem_stage(30) => 
                           new_pc_value_mem_stage_i_30_port, 
                           new_pc_value_mem_stage(29) => 
                           new_pc_value_mem_stage_i_29_port, 
                           new_pc_value_mem_stage(28) => 
                           new_pc_value_mem_stage_i_28_port, 
                           new_pc_value_mem_stage(27) => 
                           new_pc_value_mem_stage_i_27_port, 
                           new_pc_value_mem_stage(26) => 
                           new_pc_value_mem_stage_i_26_port, 
                           new_pc_value_mem_stage(25) => 
                           new_pc_value_mem_stage_i_25_port, 
                           new_pc_value_mem_stage(24) => 
                           new_pc_value_mem_stage_i_24_port, 
                           new_pc_value_mem_stage(23) => 
                           new_pc_value_mem_stage_i_23_port, 
                           new_pc_value_mem_stage(22) => 
                           new_pc_value_mem_stage_i_22_port, 
                           new_pc_value_mem_stage(21) => 
                           new_pc_value_mem_stage_i_21_port, 
                           new_pc_value_mem_stage(20) => 
                           new_pc_value_mem_stage_i_20_port, 
                           new_pc_value_mem_stage(19) => 
                           new_pc_value_mem_stage_i_19_port, 
                           new_pc_value_mem_stage(18) => 
                           new_pc_value_mem_stage_i_18_port, 
                           new_pc_value_mem_stage(17) => 
                           new_pc_value_mem_stage_i_17_port, 
                           new_pc_value_mem_stage(16) => 
                           new_pc_value_mem_stage_i_16_port, 
                           new_pc_value_mem_stage(15) => 
                           new_pc_value_mem_stage_i_15_port, 
                           new_pc_value_mem_stage(14) => 
                           new_pc_value_mem_stage_i_14_port, 
                           new_pc_value_mem_stage(13) => 
                           new_pc_value_mem_stage_i_13_port, 
                           new_pc_value_mem_stage(12) => 
                           new_pc_value_mem_stage_i_12_port, 
                           new_pc_value_mem_stage(11) => 
                           new_pc_value_mem_stage_i_11_port, 
                           new_pc_value_mem_stage(10) => 
                           new_pc_value_mem_stage_i_10_port, 
                           new_pc_value_mem_stage(9) => 
                           new_pc_value_mem_stage_i_9_port, 
                           new_pc_value_mem_stage(8) => 
                           new_pc_value_mem_stage_i_8_port, 
                           new_pc_value_mem_stage(7) => 
                           new_pc_value_mem_stage_i_7_port, 
                           new_pc_value_mem_stage(6) => 
                           new_pc_value_mem_stage_i_6_port, 
                           new_pc_value_mem_stage(5) => 
                           new_pc_value_mem_stage_i_5_port, 
                           new_pc_value_mem_stage(4) => 
                           new_pc_value_mem_stage_i_4_port, 
                           new_pc_value_mem_stage(3) => 
                           new_pc_value_mem_stage_i_3_port, 
                           new_pc_value_mem_stage(2) => 
                           new_pc_value_mem_stage_i_2_port, 
                           new_pc_value_mem_stage(1) => 
                           new_pc_value_mem_stage_i_1_port, 
                           new_pc_value_mem_stage(0) => 
                           new_pc_value_mem_stage_i_0_port, branch_taken => 
                           branch_condition_i_0_port, new_pc_value(31) => 
                           new_pc_value_decode_31_port, new_pc_value(30) => 
                           new_pc_value_decode_30_port, new_pc_value(29) => 
                           new_pc_value_decode_29_port, new_pc_value(28) => 
                           new_pc_value_decode_28_port, new_pc_value(27) => 
                           new_pc_value_decode_27_port, new_pc_value(26) => 
                           new_pc_value_decode_26_port, new_pc_value(25) => 
                           new_pc_value_decode_25_port, new_pc_value(24) => 
                           new_pc_value_decode_24_port, new_pc_value(23) => 
                           new_pc_value_decode_23_port, new_pc_value(22) => 
                           new_pc_value_decode_22_port, new_pc_value(21) => 
                           new_pc_value_decode_21_port, new_pc_value(20) => 
                           new_pc_value_decode_20_port, new_pc_value(19) => 
                           new_pc_value_decode_19_port, new_pc_value(18) => 
                           new_pc_value_decode_18_port, new_pc_value(17) => 
                           new_pc_value_decode_17_port, new_pc_value(16) => 
                           new_pc_value_decode_16_port, new_pc_value(15) => 
                           new_pc_value_decode_15_port, new_pc_value(14) => 
                           new_pc_value_decode_14_port, new_pc_value(13) => 
                           new_pc_value_decode_13_port, new_pc_value(12) => 
                           new_pc_value_decode_12_port, new_pc_value(11) => 
                           new_pc_value_decode_11_port, new_pc_value(10) => 
                           new_pc_value_decode_10_port, new_pc_value(9) => 
                           new_pc_value_decode_9_port, new_pc_value(8) => 
                           new_pc_value_decode_8_port, new_pc_value(7) => 
                           new_pc_value_decode_7_port, new_pc_value(6) => 
                           new_pc_value_decode_6_port, new_pc_value(5) => 
                           new_pc_value_decode_5_port, new_pc_value(4) => 
                           new_pc_value_decode_4_port, new_pc_value(3) => 
                           new_pc_value_decode_3_port, new_pc_value(2) => 
                           new_pc_value_decode_2_port, new_pc_value(1) => 
                           new_pc_value_decode_1_port, new_pc_value(0) => 
                           new_pc_value_decode_0_port, IRAM_ADDRESS(31) => 
                           IRAM_ADDRESS(31), IRAM_ADDRESS(30) => 
                           IRAM_ADDRESS(30), IRAM_ADDRESS(29) => 
                           IRAM_ADDRESS(29), IRAM_ADDRESS(28) => 
                           IRAM_ADDRESS(28), IRAM_ADDRESS(27) => 
                           IRAM_ADDRESS(27), IRAM_ADDRESS(26) => 
                           IRAM_ADDRESS(26), IRAM_ADDRESS(25) => 
                           IRAM_ADDRESS(25), IRAM_ADDRESS(24) => 
                           IRAM_ADDRESS(24), IRAM_ADDRESS(23) => 
                           IRAM_ADDRESS(23), IRAM_ADDRESS(22) => 
                           IRAM_ADDRESS(22), IRAM_ADDRESS(21) => 
                           IRAM_ADDRESS(21), IRAM_ADDRESS(20) => 
                           IRAM_ADDRESS(20), IRAM_ADDRESS(19) => 
                           IRAM_ADDRESS(19), IRAM_ADDRESS(18) => 
                           IRAM_ADDRESS(18), IRAM_ADDRESS(17) => 
                           IRAM_ADDRESS(17), IRAM_ADDRESS(16) => 
                           IRAM_ADDRESS(16), IRAM_ADDRESS(15) => 
                           IRAM_ADDRESS(15), IRAM_ADDRESS(14) => 
                           IRAM_ADDRESS(14), IRAM_ADDRESS(13) => 
                           IRAM_ADDRESS(13), IRAM_ADDRESS(12) => 
                           IRAM_ADDRESS(12), IRAM_ADDRESS(11) => 
                           IRAM_ADDRESS(11), IRAM_ADDRESS(10) => 
                           IRAM_ADDRESS(10), IRAM_ADDRESS(9) => IRAM_ADDRESS(9)
                           , IRAM_ADDRESS(8) => IRAM_ADDRESS(8), 
                           IRAM_ADDRESS(7) => IRAM_ADDRESS(7), IRAM_ADDRESS(6) 
                           => IRAM_ADDRESS(6), IRAM_ADDRESS(5) => 
                           IRAM_ADDRESS(5), IRAM_ADDRESS(4) => IRAM_ADDRESS(4),
                           IRAM_ADDRESS(3) => IRAM_ADDRESS(3), IRAM_ADDRESS(2) 
                           => IRAM_ADDRESS(2), IRAM_ADDRESS(1) => 
                           IRAM_ADDRESS(1), IRAM_ADDRESS(0) => IRAM_ADDRESS(0),
                           IRAM_ENABLE => IRAM_ENABLE, IRAM_READY => IRAM_READY
                           , IRAM_DATA(0) => IRAM_DATA(31), IRAM_DATA(1) => 
                           IRAM_DATA(30), IRAM_DATA(2) => IRAM_DATA(29), 
                           IRAM_DATA(3) => IRAM_DATA(28), IRAM_DATA(4) => 
                           IRAM_DATA(27), IRAM_DATA(5) => IRAM_DATA(26), 
                           IRAM_DATA(6) => IRAM_DATA(25), IRAM_DATA(7) => 
                           IRAM_DATA(24), IRAM_DATA(8) => IRAM_DATA(23), 
                           IRAM_DATA(9) => IRAM_DATA(22), IRAM_DATA(10) => 
                           IRAM_DATA(21), IRAM_DATA(11) => IRAM_DATA(20), 
                           IRAM_DATA(12) => IRAM_DATA(19), IRAM_DATA(13) => 
                           IRAM_DATA(18), IRAM_DATA(14) => IRAM_DATA(17), 
                           IRAM_DATA(15) => IRAM_DATA(16), IRAM_DATA(16) => 
                           IRAM_DATA(15), IRAM_DATA(17) => IRAM_DATA(14), 
                           IRAM_DATA(18) => IRAM_DATA(13), IRAM_DATA(19) => 
                           IRAM_DATA(12), IRAM_DATA(20) => IRAM_DATA(11), 
                           IRAM_DATA(21) => IRAM_DATA(10), IRAM_DATA(22) => 
                           IRAM_DATA(9), IRAM_DATA(23) => IRAM_DATA(8), 
                           IRAM_DATA(24) => IRAM_DATA(7), IRAM_DATA(25) => 
                           IRAM_DATA(6), IRAM_DATA(26) => IRAM_DATA(5), 
                           IRAM_DATA(27) => IRAM_DATA(4), IRAM_DATA(28) => 
                           IRAM_DATA(3), IRAM_DATA(29) => IRAM_DATA(2), 
                           IRAM_DATA(30) => IRAM_DATA(1), IRAM_DATA(31) => 
                           IRAM_DATA(0), curr_instruction(31) => 
                           curr_instruction_to_cu_31_port, curr_instruction(30)
                           => curr_instruction_to_cu_30_port, 
                           curr_instruction(29) => 
                           curr_instruction_to_cu_29_port, curr_instruction(28)
                           => curr_instruction_to_cu_28_port, 
                           curr_instruction(27) => 
                           curr_instruction_to_cu_27_port, curr_instruction(26)
                           => curr_instruction_to_cu_26_port, 
                           curr_instruction(25) => 
                           curr_instruction_to_cu_25_port, curr_instruction(24)
                           => curr_instruction_to_cu_24_port, 
                           curr_instruction(23) => 
                           curr_instruction_to_cu_23_port, curr_instruction(22)
                           => curr_instruction_to_cu_22_port, 
                           curr_instruction(21) => 
                           curr_instruction_to_cu_21_port, curr_instruction(20)
                           => curr_instruction_to_cu_20_port, 
                           curr_instruction(19) => 
                           curr_instruction_to_cu_19_port, curr_instruction(18)
                           => curr_instruction_to_cu_18_port, 
                           curr_instruction(17) => 
                           curr_instruction_to_cu_17_port, curr_instruction(16)
                           => curr_instruction_to_cu_16_port, 
                           curr_instruction(15) => 
                           curr_instruction_to_cu_15_port, curr_instruction(14)
                           => curr_instruction_to_cu_14_port, 
                           curr_instruction(13) => 
                           curr_instruction_to_cu_13_port, curr_instruction(12)
                           => curr_instruction_to_cu_12_port, 
                           curr_instruction(11) => 
                           curr_instruction_to_cu_11_port, curr_instruction(10)
                           => curr_instruction_to_cu_10_port, 
                           curr_instruction(9) => curr_instruction_to_cu_9_port
                           , curr_instruction(8) => 
                           curr_instruction_to_cu_8_port, curr_instruction(7) 
                           => curr_instruction_to_cu_7_port, 
                           curr_instruction(6) => curr_instruction_to_cu_6_port
                           , curr_instruction(5) => 
                           curr_instruction_to_cu_5_port, curr_instruction(4) 
                           => curr_instruction_to_cu_4_port, 
                           curr_instruction(3) => curr_instruction_to_cu_3_port
                           , curr_instruction(2) => 
                           curr_instruction_to_cu_2_port, curr_instruction(1) 
                           => curr_instruction_to_cu_1_port, 
                           curr_instruction(0) => curr_instruction_to_cu_0_port
                           , iram_enable_cu => iram_enable_cu, update_pc_branch
                           => update_pc_branch, stall => stall, iram_ready_cu 
                           => iram_ready_cu);
   decode_stage_dp : decode_stage_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 port map( 
                           clk => clk, rst => rst, new_prog_counter_val(31) => 
                           new_pc_value_decode_31_port, 
                           new_prog_counter_val(30) => 
                           new_pc_value_decode_30_port, 
                           new_prog_counter_val(29) => 
                           new_pc_value_decode_29_port, 
                           new_prog_counter_val(28) => 
                           new_pc_value_decode_28_port, 
                           new_prog_counter_val(27) => 
                           new_pc_value_decode_27_port, 
                           new_prog_counter_val(26) => 
                           new_pc_value_decode_26_port, 
                           new_prog_counter_val(25) => 
                           new_pc_value_decode_25_port, 
                           new_prog_counter_val(24) => 
                           new_pc_value_decode_24_port, 
                           new_prog_counter_val(23) => 
                           new_pc_value_decode_23_port, 
                           new_prog_counter_val(22) => 
                           new_pc_value_decode_22_port, 
                           new_prog_counter_val(21) => 
                           new_pc_value_decode_21_port, 
                           new_prog_counter_val(20) => 
                           new_pc_value_decode_20_port, 
                           new_prog_counter_val(19) => 
                           new_pc_value_decode_19_port, 
                           new_prog_counter_val(18) => 
                           new_pc_value_decode_18_port, 
                           new_prog_counter_val(17) => 
                           new_pc_value_decode_17_port, 
                           new_prog_counter_val(16) => 
                           new_pc_value_decode_16_port, 
                           new_prog_counter_val(15) => 
                           new_pc_value_decode_15_port, 
                           new_prog_counter_val(14) => 
                           new_pc_value_decode_14_port, 
                           new_prog_counter_val(13) => 
                           new_pc_value_decode_13_port, 
                           new_prog_counter_val(12) => 
                           new_pc_value_decode_12_port, 
                           new_prog_counter_val(11) => 
                           new_pc_value_decode_11_port, 
                           new_prog_counter_val(10) => 
                           new_pc_value_decode_10_port, new_prog_counter_val(9)
                           => new_pc_value_decode_9_port, 
                           new_prog_counter_val(8) => 
                           new_pc_value_decode_8_port, new_prog_counter_val(7) 
                           => new_pc_value_decode_7_port, 
                           new_prog_counter_val(6) => 
                           new_pc_value_decode_6_port, new_prog_counter_val(5) 
                           => new_pc_value_decode_5_port, 
                           new_prog_counter_val(4) => 
                           new_pc_value_decode_4_port, new_prog_counter_val(3) 
                           => new_pc_value_decode_3_port, 
                           new_prog_counter_val(2) => 
                           new_pc_value_decode_2_port, new_prog_counter_val(1) 
                           => new_pc_value_decode_1_port, 
                           new_prog_counter_val(0) => 
                           new_pc_value_decode_0_port, instruction_reg(31) => 
                           curr_instruction_to_cu_31_port, instruction_reg(30) 
                           => curr_instruction_to_cu_30_port, 
                           instruction_reg(29) => 
                           curr_instruction_to_cu_29_port, instruction_reg(28) 
                           => curr_instruction_to_cu_28_port, 
                           instruction_reg(27) => 
                           curr_instruction_to_cu_27_port, instruction_reg(26) 
                           => curr_instruction_to_cu_26_port, 
                           instruction_reg(25) => 
                           curr_instruction_to_cu_25_port, instruction_reg(24) 
                           => curr_instruction_to_cu_24_port, 
                           instruction_reg(23) => 
                           curr_instruction_to_cu_23_port, instruction_reg(22) 
                           => curr_instruction_to_cu_22_port, 
                           instruction_reg(21) => 
                           curr_instruction_to_cu_21_port, instruction_reg(20) 
                           => curr_instruction_to_cu_20_port, 
                           instruction_reg(19) => 
                           curr_instruction_to_cu_19_port, instruction_reg(18) 
                           => curr_instruction_to_cu_18_port, 
                           instruction_reg(17) => 
                           curr_instruction_to_cu_17_port, instruction_reg(16) 
                           => curr_instruction_to_cu_16_port, 
                           instruction_reg(15) => 
                           curr_instruction_to_cu_15_port, instruction_reg(14) 
                           => curr_instruction_to_cu_14_port, 
                           instruction_reg(13) => 
                           curr_instruction_to_cu_13_port, instruction_reg(12) 
                           => curr_instruction_to_cu_12_port, 
                           instruction_reg(11) => 
                           curr_instruction_to_cu_11_port, instruction_reg(10) 
                           => curr_instruction_to_cu_10_port, 
                           instruction_reg(9) => curr_instruction_to_cu_9_port,
                           instruction_reg(8) => curr_instruction_to_cu_8_port,
                           instruction_reg(7) => curr_instruction_to_cu_7_port,
                           instruction_reg(6) => curr_instruction_to_cu_6_port,
                           instruction_reg(5) => curr_instruction_to_cu_5_port,
                           instruction_reg(4) => curr_instruction_to_cu_4_port,
                           instruction_reg(3) => curr_instruction_to_cu_3_port,
                           instruction_reg(2) => curr_instruction_to_cu_2_port,
                           instruction_reg(1) => curr_instruction_to_cu_1_port,
                           instruction_reg(0) => curr_instruction_to_cu_0_port,
                           val_a(31) => val_a_i_31_port, val_a(30) => 
                           val_a_i_30_port, val_a(29) => val_a_i_29_port, 
                           val_a(28) => val_a_i_28_port, val_a(27) => 
                           val_a_i_27_port, val_a(26) => val_a_i_26_port, 
                           val_a(25) => val_a_i_25_port, val_a(24) => 
                           val_a_i_24_port, val_a(23) => val_a_i_23_port, 
                           val_a(22) => val_a_i_22_port, val_a(21) => 
                           val_a_i_21_port, val_a(20) => val_a_i_20_port, 
                           val_a(19) => val_a_i_19_port, val_a(18) => 
                           val_a_i_18_port, val_a(17) => val_a_i_17_port, 
                           val_a(16) => val_a_i_16_port, val_a(15) => 
                           val_a_i_15_port, val_a(14) => val_a_i_14_port, 
                           val_a(13) => val_a_i_13_port, val_a(12) => 
                           val_a_i_12_port, val_a(11) => val_a_i_11_port, 
                           val_a(10) => val_a_i_10_port, val_a(9) => 
                           val_a_i_9_port, val_a(8) => val_a_i_8_port, val_a(7)
                           => val_a_i_7_port, val_a(6) => val_a_i_6_port, 
                           val_a(5) => val_a_i_5_port, val_a(4) => 
                           val_a_i_4_port, val_a(3) => val_a_i_3_port, val_a(2)
                           => val_a_i_2_port, val_a(1) => val_a_i_1_port, 
                           val_a(0) => val_a_i_0_port, 
                           new_prog_counter_val_exe(31) => 
                           new_prog_counter_val_exe_i_31_port, 
                           new_prog_counter_val_exe(30) => 
                           new_prog_counter_val_exe_i_30_port, 
                           new_prog_counter_val_exe(29) => 
                           new_prog_counter_val_exe_i_29_port, 
                           new_prog_counter_val_exe(28) => 
                           new_prog_counter_val_exe_i_28_port, 
                           new_prog_counter_val_exe(27) => 
                           new_prog_counter_val_exe_i_27_port, 
                           new_prog_counter_val_exe(26) => 
                           new_prog_counter_val_exe_i_26_port, 
                           new_prog_counter_val_exe(25) => 
                           new_prog_counter_val_exe_i_25_port, 
                           new_prog_counter_val_exe(24) => 
                           new_prog_counter_val_exe_i_24_port, 
                           new_prog_counter_val_exe(23) => 
                           new_prog_counter_val_exe_i_23_port, 
                           new_prog_counter_val_exe(22) => 
                           new_prog_counter_val_exe_i_22_port, 
                           new_prog_counter_val_exe(21) => 
                           new_prog_counter_val_exe_i_21_port, 
                           new_prog_counter_val_exe(20) => 
                           new_prog_counter_val_exe_i_20_port, 
                           new_prog_counter_val_exe(19) => 
                           new_prog_counter_val_exe_i_19_port, 
                           new_prog_counter_val_exe(18) => 
                           new_prog_counter_val_exe_i_18_port, 
                           new_prog_counter_val_exe(17) => 
                           new_prog_counter_val_exe_i_17_port, 
                           new_prog_counter_val_exe(16) => 
                           new_prog_counter_val_exe_i_16_port, 
                           new_prog_counter_val_exe(15) => 
                           new_prog_counter_val_exe_i_15_port, 
                           new_prog_counter_val_exe(14) => 
                           new_prog_counter_val_exe_i_14_port, 
                           new_prog_counter_val_exe(13) => 
                           new_prog_counter_val_exe_i_13_port, 
                           new_prog_counter_val_exe(12) => 
                           new_prog_counter_val_exe_i_12_port, 
                           new_prog_counter_val_exe(11) => 
                           new_prog_counter_val_exe_i_11_port, 
                           new_prog_counter_val_exe(10) => 
                           new_prog_counter_val_exe_i_10_port, 
                           new_prog_counter_val_exe(9) => 
                           new_prog_counter_val_exe_i_9_port, 
                           new_prog_counter_val_exe(8) => 
                           new_prog_counter_val_exe_i_8_port, 
                           new_prog_counter_val_exe(7) => 
                           new_prog_counter_val_exe_i_7_port, 
                           new_prog_counter_val_exe(6) => 
                           new_prog_counter_val_exe_i_6_port, 
                           new_prog_counter_val_exe(5) => 
                           new_prog_counter_val_exe_i_5_port, 
                           new_prog_counter_val_exe(4) => 
                           new_prog_counter_val_exe_i_4_port, 
                           new_prog_counter_val_exe(3) => 
                           new_prog_counter_val_exe_i_3_port, 
                           new_prog_counter_val_exe(2) => 
                           new_prog_counter_val_exe_i_2_port, 
                           new_prog_counter_val_exe(1) => 
                           new_prog_counter_val_exe_i_1_port, 
                           new_prog_counter_val_exe(0) => 
                           new_prog_counter_val_exe_i_0_port, val_b(31) => 
                           val_b_i_31_port, val_b(30) => val_b_i_30_port, 
                           val_b(29) => val_b_i_29_port, val_b(28) => 
                           val_b_i_28_port, val_b(27) => val_b_i_27_port, 
                           val_b(26) => val_b_i_26_port, val_b(25) => 
                           val_b_i_25_port, val_b(24) => val_b_i_24_port, 
                           val_b(23) => val_b_i_23_port, val_b(22) => 
                           val_b_i_22_port, val_b(21) => val_b_i_21_port, 
                           val_b(20) => val_b_i_20_port, val_b(19) => 
                           val_b_i_19_port, val_b(18) => val_b_i_18_port, 
                           val_b(17) => val_b_i_17_port, val_b(16) => 
                           val_b_i_16_port, val_b(15) => val_b_i_15_port, 
                           val_b(14) => val_b_i_14_port, val_b(13) => 
                           val_b_i_13_port, val_b(12) => val_b_i_12_port, 
                           val_b(11) => val_b_i_11_port, val_b(10) => 
                           val_b_i_10_port, val_b(9) => val_b_i_9_port, 
                           val_b(8) => val_b_i_8_port, val_b(7) => 
                           val_b_i_7_port, val_b(6) => val_b_i_6_port, val_b(5)
                           => val_b_i_5_port, val_b(4) => val_b_i_4_port, 
                           val_b(3) => val_b_i_3_port, val_b(2) => 
                           val_b_i_2_port, val_b(1) => val_b_i_1_port, val_b(0)
                           => val_b_i_0_port, val_immediate(31) => 
                           val_immediate_i_31_port, val_immediate(30) => 
                           val_immediate_i_30_port, val_immediate(29) => 
                           val_immediate_i_29_port, val_immediate(28) => 
                           val_immediate_i_28_port, val_immediate(27) => 
                           val_immediate_i_27_port, val_immediate(26) => 
                           val_immediate_i_26_port, val_immediate(25) => 
                           val_immediate_i_25_port, val_immediate(24) => 
                           val_immediate_i_24_port, val_immediate(23) => 
                           val_immediate_i_23_port, val_immediate(22) => 
                           val_immediate_i_22_port, val_immediate(21) => 
                           val_immediate_i_21_port, val_immediate(20) => 
                           val_immediate_i_20_port, val_immediate(19) => 
                           val_immediate_i_19_port, val_immediate(18) => 
                           val_immediate_i_18_port, val_immediate(17) => 
                           val_immediate_i_17_port, val_immediate(16) => 
                           val_immediate_i_16_port, val_immediate(15) => 
                           val_immediate_i_15_port, val_immediate(14) => 
                           val_immediate_i_14_port, val_immediate(13) => 
                           val_immediate_i_13_port, val_immediate(12) => 
                           val_immediate_i_12_port, val_immediate(11) => 
                           val_immediate_i_11_port, val_immediate(10) => 
                           val_immediate_i_10_port, val_immediate(9) => 
                           val_immediate_i_9_port, val_immediate(8) => 
                           val_immediate_i_8_port, val_immediate(7) => 
                           val_immediate_i_7_port, val_immediate(6) => 
                           val_immediate_i_6_port, val_immediate(5) => 
                           val_immediate_i_5_port, val_immediate(4) => 
                           val_immediate_i_4_port, val_immediate(3) => 
                           val_immediate_i_3_port, val_immediate(2) => 
                           val_immediate_i_2_port, val_immediate(1) => 
                           val_immediate_i_1_port, val_immediate(0) => 
                           val_immediate_i_0_port, update_reg_value(31) => 
                           update_reg_value_i_31_port, update_reg_value(30) => 
                           update_reg_value_i_30_port, update_reg_value(29) => 
                           update_reg_value_i_29_port, update_reg_value(28) => 
                           update_reg_value_i_28_port, update_reg_value(27) => 
                           update_reg_value_i_27_port, update_reg_value(26) => 
                           update_reg_value_i_26_port, update_reg_value(25) => 
                           update_reg_value_i_25_port, update_reg_value(24) => 
                           update_reg_value_i_24_port, update_reg_value(23) => 
                           update_reg_value_i_23_port, update_reg_value(22) => 
                           update_reg_value_i_22_port, update_reg_value(21) => 
                           update_reg_value_i_21_port, update_reg_value(20) => 
                           update_reg_value_i_20_port, update_reg_value(19) => 
                           update_reg_value_i_19_port, update_reg_value(18) => 
                           update_reg_value_i_18_port, update_reg_value(17) => 
                           update_reg_value_i_17_port, update_reg_value(16) => 
                           update_reg_value_i_16_port, update_reg_value(15) => 
                           update_reg_value_i_15_port, update_reg_value(14) => 
                           update_reg_value_i_14_port, update_reg_value(13) => 
                           update_reg_value_i_13_port, update_reg_value(12) => 
                           update_reg_value_i_12_port, update_reg_value(11) => 
                           update_reg_value_i_11_port, update_reg_value(10) => 
                           update_reg_value_i_10_port, update_reg_value(9) => 
                           update_reg_value_i_9_port, update_reg_value(8) => 
                           update_reg_value_i_8_port, update_reg_value(7) => 
                           update_reg_value_i_7_port, update_reg_value(6) => 
                           update_reg_value_i_6_port, update_reg_value(5) => 
                           update_reg_value_i_5_port, update_reg_value(4) => 
                           update_reg_value_i_4_port, update_reg_value(3) => 
                           update_reg_value_i_3_port, update_reg_value(2) => 
                           update_reg_value_i_2_port, update_reg_value(1) => 
                           update_reg_value_i_1_port, update_reg_value(0) => 
                           update_reg_value_i_0_port, enable_rf => enable_rf, 
                           read_rf_p1 => read_rf_p1, read_rf_p2 => read_rf_p2, 
                           write_rf => write_rf, rtype_itypen => rtype_itypen, 
                           jump_sext => jump_sext, compute_sext => compute_sext
                           );
   execute_stage_dp : execute_stage_N32_PC_SIZE32 port map( clk => clk, rst => 
                           rst, val_a(31) => val_a_i_31_port, val_a(30) => 
                           val_a_i_30_port, val_a(29) => val_a_i_29_port, 
                           val_a(28) => val_a_i_28_port, val_a(27) => 
                           val_a_i_27_port, val_a(26) => val_a_i_26_port, 
                           val_a(25) => val_a_i_25_port, val_a(24) => 
                           val_a_i_24_port, val_a(23) => val_a_i_23_port, 
                           val_a(22) => val_a_i_22_port, val_a(21) => 
                           val_a_i_21_port, val_a(20) => val_a_i_20_port, 
                           val_a(19) => val_a_i_19_port, val_a(18) => 
                           val_a_i_18_port, val_a(17) => val_a_i_17_port, 
                           val_a(16) => val_a_i_16_port, val_a(15) => 
                           val_a_i_15_port, val_a(14) => val_a_i_14_port, 
                           val_a(13) => val_a_i_13_port, val_a(12) => 
                           val_a_i_12_port, val_a(11) => val_a_i_11_port, 
                           val_a(10) => val_a_i_10_port, val_a(9) => 
                           val_a_i_9_port, val_a(8) => val_a_i_8_port, val_a(7)
                           => val_a_i_7_port, val_a(6) => val_a_i_6_port, 
                           val_a(5) => val_a_i_5_port, val_a(4) => 
                           val_a_i_4_port, val_a(3) => val_a_i_3_port, val_a(2)
                           => val_a_i_2_port, val_a(1) => val_a_i_1_port, 
                           val_a(0) => val_a_i_0_port, val_b(31) => 
                           val_b_i_31_port, val_b(30) => val_b_i_30_port, 
                           val_b(29) => val_b_i_29_port, val_b(28) => 
                           val_b_i_28_port, val_b(27) => val_b_i_27_port, 
                           val_b(26) => val_b_i_26_port, val_b(25) => 
                           val_b_i_25_port, val_b(24) => val_b_i_24_port, 
                           val_b(23) => val_b_i_23_port, val_b(22) => 
                           val_b_i_22_port, val_b(21) => val_b_i_21_port, 
                           val_b(20) => val_b_i_20_port, val_b(19) => 
                           val_b_i_19_port, val_b(18) => val_b_i_18_port, 
                           val_b(17) => val_b_i_17_port, val_b(16) => 
                           val_b_i_16_port, val_b(15) => val_b_i_15_port, 
                           val_b(14) => val_b_i_14_port, val_b(13) => 
                           val_b_i_13_port, val_b(12) => val_b_i_12_port, 
                           val_b(11) => val_b_i_11_port, val_b(10) => 
                           val_b_i_10_port, val_b(9) => val_b_i_9_port, 
                           val_b(8) => val_b_i_8_port, val_b(7) => 
                           val_b_i_7_port, val_b(6) => val_b_i_6_port, val_b(5)
                           => val_b_i_5_port, val_b(4) => val_b_i_4_port, 
                           val_b(3) => val_b_i_3_port, val_b(2) => 
                           val_b_i_2_port, val_b(1) => val_b_i_1_port, val_b(0)
                           => val_b_i_0_port, val_immediate(31) => 
                           val_immediate_i_31_port, val_immediate(30) => 
                           val_immediate_i_30_port, val_immediate(29) => 
                           val_immediate_i_29_port, val_immediate(28) => 
                           val_immediate_i_28_port, val_immediate(27) => 
                           val_immediate_i_27_port, val_immediate(26) => 
                           val_immediate_i_26_port, val_immediate(25) => 
                           val_immediate_i_25_port, val_immediate(24) => 
                           val_immediate_i_24_port, val_immediate(23) => 
                           val_immediate_i_23_port, val_immediate(22) => 
                           val_immediate_i_22_port, val_immediate(21) => 
                           val_immediate_i_21_port, val_immediate(20) => 
                           val_immediate_i_20_port, val_immediate(19) => 
                           val_immediate_i_19_port, val_immediate(18) => 
                           val_immediate_i_18_port, val_immediate(17) => 
                           val_immediate_i_17_port, val_immediate(16) => 
                           val_immediate_i_16_port, val_immediate(15) => 
                           val_immediate_i_15_port, val_immediate(14) => 
                           val_immediate_i_14_port, val_immediate(13) => 
                           val_immediate_i_13_port, val_immediate(12) => 
                           val_immediate_i_12_port, val_immediate(11) => 
                           val_immediate_i_11_port, val_immediate(10) => 
                           val_immediate_i_10_port, val_immediate(9) => 
                           val_immediate_i_9_port, val_immediate(8) => 
                           val_immediate_i_8_port, val_immediate(7) => 
                           val_immediate_i_7_port, val_immediate(6) => 
                           val_immediate_i_6_port, val_immediate(5) => 
                           val_immediate_i_5_port, val_immediate(4) => 
                           val_immediate_i_4_port, val_immediate(3) => 
                           val_immediate_i_3_port, val_immediate(2) => 
                           val_immediate_i_2_port, val_immediate(1) => 
                           val_immediate_i_1_port, val_immediate(0) => 
                           val_immediate_i_0_port, new_prog_counter_val_exe(31)
                           => new_prog_counter_val_exe_i_31_port, 
                           new_prog_counter_val_exe(30) => 
                           new_prog_counter_val_exe_i_30_port, 
                           new_prog_counter_val_exe(29) => 
                           new_prog_counter_val_exe_i_29_port, 
                           new_prog_counter_val_exe(28) => 
                           new_prog_counter_val_exe_i_28_port, 
                           new_prog_counter_val_exe(27) => 
                           new_prog_counter_val_exe_i_27_port, 
                           new_prog_counter_val_exe(26) => 
                           new_prog_counter_val_exe_i_26_port, 
                           new_prog_counter_val_exe(25) => 
                           new_prog_counter_val_exe_i_25_port, 
                           new_prog_counter_val_exe(24) => 
                           new_prog_counter_val_exe_i_24_port, 
                           new_prog_counter_val_exe(23) => 
                           new_prog_counter_val_exe_i_23_port, 
                           new_prog_counter_val_exe(22) => 
                           new_prog_counter_val_exe_i_22_port, 
                           new_prog_counter_val_exe(21) => 
                           new_prog_counter_val_exe_i_21_port, 
                           new_prog_counter_val_exe(20) => 
                           new_prog_counter_val_exe_i_20_port, 
                           new_prog_counter_val_exe(19) => 
                           new_prog_counter_val_exe_i_19_port, 
                           new_prog_counter_val_exe(18) => 
                           new_prog_counter_val_exe_i_18_port, 
                           new_prog_counter_val_exe(17) => 
                           new_prog_counter_val_exe_i_17_port, 
                           new_prog_counter_val_exe(16) => 
                           new_prog_counter_val_exe_i_16_port, 
                           new_prog_counter_val_exe(15) => 
                           new_prog_counter_val_exe_i_15_port, 
                           new_prog_counter_val_exe(14) => 
                           new_prog_counter_val_exe_i_14_port, 
                           new_prog_counter_val_exe(13) => 
                           new_prog_counter_val_exe_i_13_port, 
                           new_prog_counter_val_exe(12) => 
                           new_prog_counter_val_exe_i_12_port, 
                           new_prog_counter_val_exe(11) => 
                           new_prog_counter_val_exe_i_11_port, 
                           new_prog_counter_val_exe(10) => 
                           new_prog_counter_val_exe_i_10_port, 
                           new_prog_counter_val_exe(9) => 
                           new_prog_counter_val_exe_i_9_port, 
                           new_prog_counter_val_exe(8) => 
                           new_prog_counter_val_exe_i_8_port, 
                           new_prog_counter_val_exe(7) => 
                           new_prog_counter_val_exe_i_7_port, 
                           new_prog_counter_val_exe(6) => 
                           new_prog_counter_val_exe_i_6_port, 
                           new_prog_counter_val_exe(5) => 
                           new_prog_counter_val_exe_i_5_port, 
                           new_prog_counter_val_exe(4) => 
                           new_prog_counter_val_exe_i_4_port, 
                           new_prog_counter_val_exe(3) => 
                           new_prog_counter_val_exe_i_3_port, 
                           new_prog_counter_val_exe(2) => 
                           new_prog_counter_val_exe_i_2_port, 
                           new_prog_counter_val_exe(1) => 
                           new_prog_counter_val_exe_i_1_port, 
                           new_prog_counter_val_exe(0) => 
                           new_prog_counter_val_exe_i_0_port, branch_condition 
                           => branch_condition_i_0_port, 
                           prog_counter_forwaded(31) => 
                           prog_counter_forwaded_i_31_port, 
                           prog_counter_forwaded(30) => 
                           prog_counter_forwaded_i_30_port, 
                           prog_counter_forwaded(29) => 
                           prog_counter_forwaded_i_29_port, 
                           prog_counter_forwaded(28) => 
                           prog_counter_forwaded_i_28_port, 
                           prog_counter_forwaded(27) => 
                           prog_counter_forwaded_i_27_port, 
                           prog_counter_forwaded(26) => 
                           prog_counter_forwaded_i_26_port, 
                           prog_counter_forwaded(25) => 
                           prog_counter_forwaded_i_25_port, 
                           prog_counter_forwaded(24) => 
                           prog_counter_forwaded_i_24_port, 
                           prog_counter_forwaded(23) => 
                           prog_counter_forwaded_i_23_port, 
                           prog_counter_forwaded(22) => 
                           prog_counter_forwaded_i_22_port, 
                           prog_counter_forwaded(21) => 
                           prog_counter_forwaded_i_21_port, 
                           prog_counter_forwaded(20) => 
                           prog_counter_forwaded_i_20_port, 
                           prog_counter_forwaded(19) => 
                           prog_counter_forwaded_i_19_port, 
                           prog_counter_forwaded(18) => 
                           prog_counter_forwaded_i_18_port, 
                           prog_counter_forwaded(17) => 
                           prog_counter_forwaded_i_17_port, 
                           prog_counter_forwaded(16) => 
                           prog_counter_forwaded_i_16_port, 
                           prog_counter_forwaded(15) => 
                           prog_counter_forwaded_i_15_port, 
                           prog_counter_forwaded(14) => 
                           prog_counter_forwaded_i_14_port, 
                           prog_counter_forwaded(13) => 
                           prog_counter_forwaded_i_13_port, 
                           prog_counter_forwaded(12) => 
                           prog_counter_forwaded_i_12_port, 
                           prog_counter_forwaded(11) => 
                           prog_counter_forwaded_i_11_port, 
                           prog_counter_forwaded(10) => 
                           prog_counter_forwaded_i_10_port, 
                           prog_counter_forwaded(9) => 
                           prog_counter_forwaded_i_9_port, 
                           prog_counter_forwaded(8) => 
                           prog_counter_forwaded_i_8_port, 
                           prog_counter_forwaded(7) => 
                           prog_counter_forwaded_i_7_port, 
                           prog_counter_forwaded(6) => 
                           prog_counter_forwaded_i_6_port, 
                           prog_counter_forwaded(5) => 
                           prog_counter_forwaded_i_5_port, 
                           prog_counter_forwaded(4) => 
                           prog_counter_forwaded_i_4_port, 
                           prog_counter_forwaded(3) => 
                           prog_counter_forwaded_i_3_port, 
                           prog_counter_forwaded(2) => 
                           prog_counter_forwaded_i_2_port, 
                           prog_counter_forwaded(1) => 
                           prog_counter_forwaded_i_1_port, 
                           prog_counter_forwaded(0) => 
                           prog_counter_forwaded_i_0_port, alu_output_val(31) 
                           => alu_output_val_i_31_port, alu_output_val(30) => 
                           alu_output_val_i_30_port, alu_output_val(29) => 
                           alu_output_val_i_29_port, alu_output_val(28) => 
                           alu_output_val_i_28_port, alu_output_val(27) => 
                           alu_output_val_i_27_port, alu_output_val(26) => 
                           alu_output_val_i_26_port, alu_output_val(25) => 
                           alu_output_val_i_25_port, alu_output_val(24) => 
                           alu_output_val_i_24_port, alu_output_val(23) => 
                           alu_output_val_i_23_port, alu_output_val(22) => 
                           alu_output_val_i_22_port, alu_output_val(21) => 
                           alu_output_val_i_21_port, alu_output_val(20) => 
                           alu_output_val_i_20_port, alu_output_val(19) => 
                           alu_output_val_i_19_port, alu_output_val(18) => 
                           alu_output_val_i_18_port, alu_output_val(17) => 
                           alu_output_val_i_17_port, alu_output_val(16) => 
                           alu_output_val_i_16_port, alu_output_val(15) => 
                           alu_output_val_i_15_port, alu_output_val(14) => 
                           alu_output_val_i_14_port, alu_output_val(13) => 
                           alu_output_val_i_13_port, alu_output_val(12) => 
                           alu_output_val_i_12_port, alu_output_val(11) => 
                           alu_output_val_i_11_port, alu_output_val(10) => 
                           alu_output_val_i_10_port, alu_output_val(9) => 
                           alu_output_val_i_9_port, alu_output_val(8) => 
                           alu_output_val_i_8_port, alu_output_val(7) => 
                           alu_output_val_i_7_port, alu_output_val(6) => 
                           alu_output_val_i_6_port, alu_output_val(5) => 
                           alu_output_val_i_5_port, alu_output_val(4) => 
                           alu_output_val_i_4_port, alu_output_val(3) => 
                           alu_output_val_i_3_port, alu_output_val(2) => 
                           alu_output_val_i_2_port, alu_output_val(1) => 
                           alu_output_val_i_1_port, alu_output_val(0) => 
                           alu_output_val_i_0_port, value_to_mem(31) => 
                           value_to_mem_i_31_port, value_to_mem(30) => 
                           value_to_mem_i_30_port, value_to_mem(29) => 
                           value_to_mem_i_29_port, value_to_mem(28) => 
                           value_to_mem_i_28_port, value_to_mem(27) => 
                           value_to_mem_i_27_port, value_to_mem(26) => 
                           value_to_mem_i_26_port, value_to_mem(25) => 
                           value_to_mem_i_25_port, value_to_mem(24) => 
                           value_to_mem_i_24_port, value_to_mem(23) => 
                           value_to_mem_i_23_port, value_to_mem(22) => 
                           value_to_mem_i_22_port, value_to_mem(21) => 
                           value_to_mem_i_21_port, value_to_mem(20) => 
                           value_to_mem_i_20_port, value_to_mem(19) => 
                           value_to_mem_i_19_port, value_to_mem(18) => 
                           value_to_mem_i_18_port, value_to_mem(17) => 
                           value_to_mem_i_17_port, value_to_mem(16) => 
                           value_to_mem_i_16_port, value_to_mem(15) => 
                           value_to_mem_i_15_port, value_to_mem(14) => 
                           value_to_mem_i_14_port, value_to_mem(13) => 
                           value_to_mem_i_13_port, value_to_mem(12) => 
                           value_to_mem_i_12_port, value_to_mem(11) => 
                           value_to_mem_i_11_port, value_to_mem(10) => 
                           value_to_mem_i_10_port, value_to_mem(9) => 
                           value_to_mem_i_9_port, value_to_mem(8) => 
                           value_to_mem_i_8_port, value_to_mem(7) => 
                           value_to_mem_i_7_port, value_to_mem(6) => 
                           value_to_mem_i_6_port, value_to_mem(5) => 
                           value_to_mem_i_5_port, value_to_mem(4) => 
                           value_to_mem_i_4_port, value_to_mem(3) => 
                           value_to_mem_i_3_port, value_to_mem(2) => 
                           value_to_mem_i_2_port, value_to_mem(1) => 
                           value_to_mem_i_1_port, value_to_mem(0) => 
                           value_to_mem_i_0_port, signed_notsigned => 
                           signed_notsigned, alu_op_type(3) => alu_op_type(3), 
                           alu_op_type(2) => alu_op_type(2), alu_op_type(1) => 
                           alu_op_type(1), alu_op_type(0) => alu_op_type(0), 
                           sel_val_a => sel_val_a, sel_val_b => sel_val_b, cin 
                           => alu_cin, overflow => alu_overflow, 
                           zero_mul_detect => zero_mul_detect, mul_exeception 
                           => mul_exeception, evaluate_branch(1) => 
                           evaluate_branch(1), evaluate_branch(0) => 
                           evaluate_branch(0));
   memory_stage_dp : memory_stage_N32_PC_SIZE32 port map( clk => clk, rst => 
                           rst, new_pc_value(31) => 
                           prog_counter_forwaded_i_31_port, new_pc_value(30) =>
                           prog_counter_forwaded_i_30_port, new_pc_value(29) =>
                           prog_counter_forwaded_i_29_port, new_pc_value(28) =>
                           prog_counter_forwaded_i_28_port, new_pc_value(27) =>
                           prog_counter_forwaded_i_27_port, new_pc_value(26) =>
                           prog_counter_forwaded_i_26_port, new_pc_value(25) =>
                           prog_counter_forwaded_i_25_port, new_pc_value(24) =>
                           prog_counter_forwaded_i_24_port, new_pc_value(23) =>
                           prog_counter_forwaded_i_23_port, new_pc_value(22) =>
                           prog_counter_forwaded_i_22_port, new_pc_value(21) =>
                           prog_counter_forwaded_i_21_port, new_pc_value(20) =>
                           prog_counter_forwaded_i_20_port, new_pc_value(19) =>
                           prog_counter_forwaded_i_19_port, new_pc_value(18) =>
                           prog_counter_forwaded_i_18_port, new_pc_value(17) =>
                           prog_counter_forwaded_i_17_port, new_pc_value(16) =>
                           prog_counter_forwaded_i_16_port, new_pc_value(15) =>
                           prog_counter_forwaded_i_15_port, new_pc_value(14) =>
                           prog_counter_forwaded_i_14_port, new_pc_value(13) =>
                           prog_counter_forwaded_i_13_port, new_pc_value(12) =>
                           prog_counter_forwaded_i_12_port, new_pc_value(11) =>
                           prog_counter_forwaded_i_11_port, new_pc_value(10) =>
                           prog_counter_forwaded_i_10_port, new_pc_value(9) => 
                           prog_counter_forwaded_i_9_port, new_pc_value(8) => 
                           prog_counter_forwaded_i_8_port, new_pc_value(7) => 
                           prog_counter_forwaded_i_7_port, new_pc_value(6) => 
                           prog_counter_forwaded_i_6_port, new_pc_value(5) => 
                           prog_counter_forwaded_i_5_port, new_pc_value(4) => 
                           prog_counter_forwaded_i_4_port, new_pc_value(3) => 
                           prog_counter_forwaded_i_3_port, new_pc_value(2) => 
                           prog_counter_forwaded_i_2_port, new_pc_value(1) => 
                           prog_counter_forwaded_i_1_port, new_pc_value(0) => 
                           prog_counter_forwaded_i_0_port, 
                           new_pc_value_branch(31) => 
                           new_pc_value_mem_stage_i_31_port, 
                           new_pc_value_branch(30) => 
                           new_pc_value_mem_stage_i_30_port, 
                           new_pc_value_branch(29) => 
                           new_pc_value_mem_stage_i_29_port, 
                           new_pc_value_branch(28) => 
                           new_pc_value_mem_stage_i_28_port, 
                           new_pc_value_branch(27) => 
                           new_pc_value_mem_stage_i_27_port, 
                           new_pc_value_branch(26) => 
                           new_pc_value_mem_stage_i_26_port, 
                           new_pc_value_branch(25) => 
                           new_pc_value_mem_stage_i_25_port, 
                           new_pc_value_branch(24) => 
                           new_pc_value_mem_stage_i_24_port, 
                           new_pc_value_branch(23) => 
                           new_pc_value_mem_stage_i_23_port, 
                           new_pc_value_branch(22) => 
                           new_pc_value_mem_stage_i_22_port, 
                           new_pc_value_branch(21) => 
                           new_pc_value_mem_stage_i_21_port, 
                           new_pc_value_branch(20) => 
                           new_pc_value_mem_stage_i_20_port, 
                           new_pc_value_branch(19) => 
                           new_pc_value_mem_stage_i_19_port, 
                           new_pc_value_branch(18) => 
                           new_pc_value_mem_stage_i_18_port, 
                           new_pc_value_branch(17) => 
                           new_pc_value_mem_stage_i_17_port, 
                           new_pc_value_branch(16) => 
                           new_pc_value_mem_stage_i_16_port, 
                           new_pc_value_branch(15) => 
                           new_pc_value_mem_stage_i_15_port, 
                           new_pc_value_branch(14) => 
                           new_pc_value_mem_stage_i_14_port, 
                           new_pc_value_branch(13) => 
                           new_pc_value_mem_stage_i_13_port, 
                           new_pc_value_branch(12) => 
                           new_pc_value_mem_stage_i_12_port, 
                           new_pc_value_branch(11) => 
                           new_pc_value_mem_stage_i_11_port, 
                           new_pc_value_branch(10) => 
                           new_pc_value_mem_stage_i_10_port, 
                           new_pc_value_branch(9) => 
                           new_pc_value_mem_stage_i_9_port, 
                           new_pc_value_branch(8) => 
                           new_pc_value_mem_stage_i_8_port, 
                           new_pc_value_branch(7) => 
                           new_pc_value_mem_stage_i_7_port, 
                           new_pc_value_branch(6) => 
                           new_pc_value_mem_stage_i_6_port, 
                           new_pc_value_branch(5) => 
                           new_pc_value_mem_stage_i_5_port, 
                           new_pc_value_branch(4) => 
                           new_pc_value_mem_stage_i_4_port, 
                           new_pc_value_branch(3) => 
                           new_pc_value_mem_stage_i_3_port, 
                           new_pc_value_branch(2) => 
                           new_pc_value_mem_stage_i_2_port, 
                           new_pc_value_branch(1) => 
                           new_pc_value_mem_stage_i_1_port, 
                           new_pc_value_branch(0) => 
                           new_pc_value_mem_stage_i_0_port, select_pc => 
                           branch_condition_i_0_port, alu_output_val(31) => 
                           alu_output_val_i_31_port, alu_output_val(30) => 
                           alu_output_val_i_30_port, alu_output_val(29) => 
                           alu_output_val_i_29_port, alu_output_val(28) => 
                           alu_output_val_i_28_port, alu_output_val(27) => 
                           alu_output_val_i_27_port, alu_output_val(26) => 
                           alu_output_val_i_26_port, alu_output_val(25) => 
                           alu_output_val_i_25_port, alu_output_val(24) => 
                           alu_output_val_i_24_port, alu_output_val(23) => 
                           alu_output_val_i_23_port, alu_output_val(22) => 
                           alu_output_val_i_22_port, alu_output_val(21) => 
                           alu_output_val_i_21_port, alu_output_val(20) => 
                           alu_output_val_i_20_port, alu_output_val(19) => 
                           alu_output_val_i_19_port, alu_output_val(18) => 
                           alu_output_val_i_18_port, alu_output_val(17) => 
                           alu_output_val_i_17_port, alu_output_val(16) => 
                           alu_output_val_i_16_port, alu_output_val(15) => 
                           alu_output_val_i_15_port, alu_output_val(14) => 
                           alu_output_val_i_14_port, alu_output_val(13) => 
                           alu_output_val_i_13_port, alu_output_val(12) => 
                           alu_output_val_i_12_port, alu_output_val(11) => 
                           alu_output_val_i_11_port, alu_output_val(10) => 
                           alu_output_val_i_10_port, alu_output_val(9) => 
                           alu_output_val_i_9_port, alu_output_val(8) => 
                           alu_output_val_i_8_port, alu_output_val(7) => 
                           alu_output_val_i_7_port, alu_output_val(6) => 
                           alu_output_val_i_6_port, alu_output_val(5) => 
                           alu_output_val_i_5_port, alu_output_val(4) => 
                           alu_output_val_i_4_port, alu_output_val(3) => 
                           alu_output_val_i_3_port, alu_output_val(2) => 
                           alu_output_val_i_2_port, alu_output_val(1) => 
                           alu_output_val_i_1_port, alu_output_val(0) => 
                           alu_output_val_i_0_port, value_to_mem(31) => 
                           value_to_mem_i_31_port, value_to_mem(30) => 
                           value_to_mem_i_30_port, value_to_mem(29) => 
                           value_to_mem_i_29_port, value_to_mem(28) => 
                           value_to_mem_i_28_port, value_to_mem(27) => 
                           value_to_mem_i_27_port, value_to_mem(26) => 
                           value_to_mem_i_26_port, value_to_mem(25) => 
                           value_to_mem_i_25_port, value_to_mem(24) => 
                           value_to_mem_i_24_port, value_to_mem(23) => 
                           value_to_mem_i_23_port, value_to_mem(22) => 
                           value_to_mem_i_22_port, value_to_mem(21) => 
                           value_to_mem_i_21_port, value_to_mem(20) => 
                           value_to_mem_i_20_port, value_to_mem(19) => 
                           value_to_mem_i_19_port, value_to_mem(18) => 
                           value_to_mem_i_18_port, value_to_mem(17) => 
                           value_to_mem_i_17_port, value_to_mem(16) => 
                           value_to_mem_i_16_port, value_to_mem(15) => 
                           value_to_mem_i_15_port, value_to_mem(14) => 
                           value_to_mem_i_14_port, value_to_mem(13) => 
                           value_to_mem_i_13_port, value_to_mem(12) => 
                           value_to_mem_i_12_port, value_to_mem(11) => 
                           value_to_mem_i_11_port, value_to_mem(10) => 
                           value_to_mem_i_10_port, value_to_mem(9) => 
                           value_to_mem_i_9_port, value_to_mem(8) => 
                           value_to_mem_i_8_port, value_to_mem(7) => 
                           value_to_mem_i_7_port, value_to_mem(6) => 
                           value_to_mem_i_6_port, value_to_mem(5) => 
                           value_to_mem_i_5_port, value_to_mem(4) => 
                           value_to_mem_i_4_port, value_to_mem(3) => 
                           value_to_mem_i_3_port, value_to_mem(2) => 
                           value_to_mem_i_2_port, value_to_mem(1) => 
                           value_to_mem_i_1_port, value_to_mem(0) => 
                           value_to_mem_i_0_port, data_from_memory(31) => 
                           data_from_memory_i_31_port, data_from_memory(30) => 
                           data_from_memory_i_30_port, data_from_memory(29) => 
                           data_from_memory_i_29_port, data_from_memory(28) => 
                           data_from_memory_i_28_port, data_from_memory(27) => 
                           data_from_memory_i_27_port, data_from_memory(26) => 
                           data_from_memory_i_26_port, data_from_memory(25) => 
                           data_from_memory_i_25_port, data_from_memory(24) => 
                           data_from_memory_i_24_port, data_from_memory(23) => 
                           data_from_memory_i_23_port, data_from_memory(22) => 
                           data_from_memory_i_22_port, data_from_memory(21) => 
                           data_from_memory_i_21_port, data_from_memory(20) => 
                           data_from_memory_i_20_port, data_from_memory(19) => 
                           data_from_memory_i_19_port, data_from_memory(18) => 
                           data_from_memory_i_18_port, data_from_memory(17) => 
                           data_from_memory_i_17_port, data_from_memory(16) => 
                           data_from_memory_i_16_port, data_from_memory(15) => 
                           data_from_memory_i_15_port, data_from_memory(14) => 
                           data_from_memory_i_14_port, data_from_memory(13) => 
                           data_from_memory_i_13_port, data_from_memory(12) => 
                           data_from_memory_i_12_port, data_from_memory(11) => 
                           data_from_memory_i_11_port, data_from_memory(10) => 
                           data_from_memory_i_10_port, data_from_memory(9) => 
                           data_from_memory_i_9_port, data_from_memory(8) => 
                           data_from_memory_i_8_port, data_from_memory(7) => 
                           data_from_memory_i_7_port, data_from_memory(6) => 
                           data_from_memory_i_6_port, data_from_memory(5) => 
                           data_from_memory_i_5_port, data_from_memory(4) => 
                           data_from_memory_i_4_port, data_from_memory(3) => 
                           data_from_memory_i_3_port, data_from_memory(2) => 
                           data_from_memory_i_2_port, data_from_memory(1) => 
                           data_from_memory_i_1_port, data_from_memory(0) => 
                           data_from_memory_i_0_port, data_from_alu(31) => 
                           data_from_alu_i_31_port, data_from_alu(30) => 
                           data_from_alu_i_30_port, data_from_alu(29) => 
                           data_from_alu_i_29_port, data_from_alu(28) => 
                           data_from_alu_i_28_port, data_from_alu(27) => 
                           data_from_alu_i_27_port, data_from_alu(26) => 
                           data_from_alu_i_26_port, data_from_alu(25) => 
                           data_from_alu_i_25_port, data_from_alu(24) => 
                           data_from_alu_i_24_port, data_from_alu(23) => 
                           data_from_alu_i_23_port, data_from_alu(22) => 
                           data_from_alu_i_22_port, data_from_alu(21) => 
                           data_from_alu_i_21_port, data_from_alu(20) => 
                           data_from_alu_i_20_port, data_from_alu(19) => 
                           data_from_alu_i_19_port, data_from_alu(18) => 
                           data_from_alu_i_18_port, data_from_alu(17) => 
                           data_from_alu_i_17_port, data_from_alu(16) => 
                           data_from_alu_i_16_port, data_from_alu(15) => 
                           data_from_alu_i_15_port, data_from_alu(14) => 
                           data_from_alu_i_14_port, data_from_alu(13) => 
                           data_from_alu_i_13_port, data_from_alu(12) => 
                           data_from_alu_i_12_port, data_from_alu(11) => 
                           data_from_alu_i_11_port, data_from_alu(10) => 
                           data_from_alu_i_10_port, data_from_alu(9) => 
                           data_from_alu_i_9_port, data_from_alu(8) => 
                           data_from_alu_i_8_port, data_from_alu(7) => 
                           data_from_alu_i_7_port, data_from_alu(6) => 
                           data_from_alu_i_6_port, data_from_alu(5) => 
                           data_from_alu_i_5_port, data_from_alu(4) => 
                           data_from_alu_i_4_port, data_from_alu(3) => 
                           data_from_alu_i_3_port, data_from_alu(2) => 
                           data_from_alu_i_2_port, data_from_alu(1) => 
                           data_from_alu_i_1_port, data_from_alu(0) => 
                           data_from_alu_i_0_port, dram_enable_cu => 
                           dram_enable_cu, dram_r_nw_cu => dram_r_nw_cu, 
                           dram_ready_cu => dram_ready_cu, DRAM_ADDRESS(31) => 
                           DRAM_ADDRESS(31), DRAM_ADDRESS(30) => 
                           DRAM_ADDRESS(30), DRAM_ADDRESS(29) => 
                           DRAM_ADDRESS(29), DRAM_ADDRESS(28) => 
                           DRAM_ADDRESS(28), DRAM_ADDRESS(27) => 
                           DRAM_ADDRESS(27), DRAM_ADDRESS(26) => 
                           DRAM_ADDRESS(26), DRAM_ADDRESS(25) => 
                           DRAM_ADDRESS(25), DRAM_ADDRESS(24) => 
                           DRAM_ADDRESS(24), DRAM_ADDRESS(23) => 
                           DRAM_ADDRESS(23), DRAM_ADDRESS(22) => 
                           DRAM_ADDRESS(22), DRAM_ADDRESS(21) => 
                           DRAM_ADDRESS(21), DRAM_ADDRESS(20) => 
                           DRAM_ADDRESS(20), DRAM_ADDRESS(19) => 
                           DRAM_ADDRESS(19), DRAM_ADDRESS(18) => 
                           DRAM_ADDRESS(18), DRAM_ADDRESS(17) => 
                           DRAM_ADDRESS(17), DRAM_ADDRESS(16) => 
                           DRAM_ADDRESS(16), DRAM_ADDRESS(15) => 
                           DRAM_ADDRESS(15), DRAM_ADDRESS(14) => 
                           DRAM_ADDRESS(14), DRAM_ADDRESS(13) => 
                           DRAM_ADDRESS(13), DRAM_ADDRESS(12) => 
                           DRAM_ADDRESS(12), DRAM_ADDRESS(11) => 
                           DRAM_ADDRESS(11), DRAM_ADDRESS(10) => 
                           DRAM_ADDRESS(10), DRAM_ADDRESS(9) => DRAM_ADDRESS(9)
                           , DRAM_ADDRESS(8) => DRAM_ADDRESS(8), 
                           DRAM_ADDRESS(7) => DRAM_ADDRESS(7), DRAM_ADDRESS(6) 
                           => DRAM_ADDRESS(6), DRAM_ADDRESS(5) => 
                           DRAM_ADDRESS(5), DRAM_ADDRESS(4) => DRAM_ADDRESS(4),
                           DRAM_ADDRESS(3) => DRAM_ADDRESS(3), DRAM_ADDRESS(2) 
                           => DRAM_ADDRESS(2), DRAM_ADDRESS(1) => n_5536, 
                           DRAM_ADDRESS(0) => n_5537, DRAM_ENABLE => 
                           DRAM_ENABLE, DRAM_READNOTWRITE => DRAM_READNOTWRITE,
                           DRAM_READY => DRAM_READY, DRAM_DATA(31) => 
                           DRAM_DATA(31), DRAM_DATA(30) => DRAM_DATA(30), 
                           DRAM_DATA(29) => DRAM_DATA(29), DRAM_DATA(28) => 
                           DRAM_DATA(28), DRAM_DATA(27) => DRAM_DATA(27), 
                           DRAM_DATA(26) => DRAM_DATA(26), DRAM_DATA(25) => 
                           DRAM_DATA(25), DRAM_DATA(24) => DRAM_DATA(24), 
                           DRAM_DATA(23) => DRAM_DATA(23), DRAM_DATA(22) => 
                           DRAM_DATA(22), DRAM_DATA(21) => DRAM_DATA(21), 
                           DRAM_DATA(20) => DRAM_DATA(20), DRAM_DATA(19) => 
                           DRAM_DATA(19), DRAM_DATA(18) => DRAM_DATA(18), 
                           DRAM_DATA(17) => DRAM_DATA(17), DRAM_DATA(16) => 
                           DRAM_DATA(16), DRAM_DATA(15) => DRAM_DATA(15), 
                           DRAM_DATA(14) => DRAM_DATA(14), DRAM_DATA(13) => 
                           DRAM_DATA(13), DRAM_DATA(12) => DRAM_DATA(12), 
                           DRAM_DATA(11) => DRAM_DATA(11), DRAM_DATA(10) => 
                           DRAM_DATA(10), DRAM_DATA(9) => DRAM_DATA(9), 
                           DRAM_DATA(8) => DRAM_DATA(8), DRAM_DATA(7) => 
                           DRAM_DATA(7), DRAM_DATA(6) => DRAM_DATA(6), 
                           DRAM_DATA(5) => DRAM_DATA(5), DRAM_DATA(4) => 
                           DRAM_DATA(4), DRAM_DATA(3) => DRAM_DATA(3), 
                           DRAM_DATA(2) => DRAM_DATA(2), DRAM_DATA(1) => 
                           DRAM_DATA(1), DRAM_DATA(0) => DRAM_DATA(0));
   write_back_stage_dp : write_back_stage_N32 port map( data_from_memory(31) =>
                           data_from_memory_i_31_port, data_from_memory(30) => 
                           data_from_memory_i_30_port, data_from_memory(29) => 
                           data_from_memory_i_29_port, data_from_memory(28) => 
                           data_from_memory_i_28_port, data_from_memory(27) => 
                           data_from_memory_i_27_port, data_from_memory(26) => 
                           data_from_memory_i_26_port, data_from_memory(25) => 
                           data_from_memory_i_25_port, data_from_memory(24) => 
                           data_from_memory_i_24_port, data_from_memory(23) => 
                           data_from_memory_i_23_port, data_from_memory(22) => 
                           data_from_memory_i_22_port, data_from_memory(21) => 
                           data_from_memory_i_21_port, data_from_memory(20) => 
                           data_from_memory_i_20_port, data_from_memory(19) => 
                           data_from_memory_i_19_port, data_from_memory(18) => 
                           data_from_memory_i_18_port, data_from_memory(17) => 
                           data_from_memory_i_17_port, data_from_memory(16) => 
                           data_from_memory_i_16_port, data_from_memory(15) => 
                           data_from_memory_i_15_port, data_from_memory(14) => 
                           data_from_memory_i_14_port, data_from_memory(13) => 
                           data_from_memory_i_13_port, data_from_memory(12) => 
                           data_from_memory_i_12_port, data_from_memory(11) => 
                           data_from_memory_i_11_port, data_from_memory(10) => 
                           data_from_memory_i_10_port, data_from_memory(9) => 
                           data_from_memory_i_9_port, data_from_memory(8) => 
                           data_from_memory_i_8_port, data_from_memory(7) => 
                           data_from_memory_i_7_port, data_from_memory(6) => 
                           data_from_memory_i_6_port, data_from_memory(5) => 
                           data_from_memory_i_5_port, data_from_memory(4) => 
                           data_from_memory_i_4_port, data_from_memory(3) => 
                           data_from_memory_i_3_port, data_from_memory(2) => 
                           data_from_memory_i_2_port, data_from_memory(1) => 
                           data_from_memory_i_1_port, data_from_memory(0) => 
                           data_from_memory_i_0_port, data_from_alu(31) => 
                           data_from_alu_i_31_port, data_from_alu(30) => 
                           data_from_alu_i_30_port, data_from_alu(29) => 
                           data_from_alu_i_29_port, data_from_alu(28) => 
                           data_from_alu_i_28_port, data_from_alu(27) => 
                           data_from_alu_i_27_port, data_from_alu(26) => 
                           data_from_alu_i_26_port, data_from_alu(25) => 
                           data_from_alu_i_25_port, data_from_alu(24) => 
                           data_from_alu_i_24_port, data_from_alu(23) => 
                           data_from_alu_i_23_port, data_from_alu(22) => 
                           data_from_alu_i_22_port, data_from_alu(21) => 
                           data_from_alu_i_21_port, data_from_alu(20) => 
                           data_from_alu_i_20_port, data_from_alu(19) => 
                           data_from_alu_i_19_port, data_from_alu(18) => 
                           data_from_alu_i_18_port, data_from_alu(17) => 
                           data_from_alu_i_17_port, data_from_alu(16) => 
                           data_from_alu_i_16_port, data_from_alu(15) => 
                           data_from_alu_i_15_port, data_from_alu(14) => 
                           data_from_alu_i_14_port, data_from_alu(13) => 
                           data_from_alu_i_13_port, data_from_alu(12) => 
                           data_from_alu_i_12_port, data_from_alu(11) => 
                           data_from_alu_i_11_port, data_from_alu(10) => 
                           data_from_alu_i_10_port, data_from_alu(9) => 
                           data_from_alu_i_9_port, data_from_alu(8) => 
                           data_from_alu_i_8_port, data_from_alu(7) => 
                           data_from_alu_i_7_port, data_from_alu(6) => 
                           data_from_alu_i_6_port, data_from_alu(5) => 
                           data_from_alu_i_5_port, data_from_alu(4) => 
                           data_from_alu_i_4_port, data_from_alu(3) => 
                           data_from_alu_i_3_port, data_from_alu(2) => 
                           data_from_alu_i_2_port, data_from_alu(1) => 
                           data_from_alu_i_1_port, data_from_alu(0) => 
                           data_from_alu_i_0_port, data_to_rf(31) => 
                           update_reg_value_i_31_port, data_to_rf(30) => 
                           update_reg_value_i_30_port, data_to_rf(29) => 
                           update_reg_value_i_29_port, data_to_rf(28) => 
                           update_reg_value_i_28_port, data_to_rf(27) => 
                           update_reg_value_i_27_port, data_to_rf(26) => 
                           update_reg_value_i_26_port, data_to_rf(25) => 
                           update_reg_value_i_25_port, data_to_rf(24) => 
                           update_reg_value_i_24_port, data_to_rf(23) => 
                           update_reg_value_i_23_port, data_to_rf(22) => 
                           update_reg_value_i_22_port, data_to_rf(21) => 
                           update_reg_value_i_21_port, data_to_rf(20) => 
                           update_reg_value_i_20_port, data_to_rf(19) => 
                           update_reg_value_i_19_port, data_to_rf(18) => 
                           update_reg_value_i_18_port, data_to_rf(17) => 
                           update_reg_value_i_17_port, data_to_rf(16) => 
                           update_reg_value_i_16_port, data_to_rf(15) => 
                           update_reg_value_i_15_port, data_to_rf(14) => 
                           update_reg_value_i_14_port, data_to_rf(13) => 
                           update_reg_value_i_13_port, data_to_rf(12) => 
                           update_reg_value_i_12_port, data_to_rf(11) => 
                           update_reg_value_i_11_port, data_to_rf(10) => 
                           update_reg_value_i_10_port, data_to_rf(9) => 
                           update_reg_value_i_9_port, data_to_rf(8) => 
                           update_reg_value_i_8_port, data_to_rf(7) => 
                           update_reg_value_i_7_port, data_to_rf(6) => 
                           update_reg_value_i_6_port, data_to_rf(5) => 
                           update_reg_value_i_5_port, data_to_rf(4) => 
                           update_reg_value_i_4_port, data_to_rf(3) => 
                           update_reg_value_i_3_port, data_to_rf(2) => 
                           update_reg_value_i_2_port, data_to_rf(1) => 
                           update_reg_value_i_1_port, data_to_rf(0) => 
                           update_reg_value_i_0_port, select_wb => select_wb);
   DRAM_ADDRESS(0) <= '0';
   DRAM_ADDRESS(1) <= '0';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity control_unit_PC_SIZE32_RF_REGS32_IR_SIZE32_CW_SIZE22 is

   port( clk, rst : in std_logic;  iram_enable_cu : out std_logic;  
         iram_ready_cu : in std_logic;  curr_instruction_to_cu : in 
         std_logic_vector (31 downto 0);  stall_pip, enable_rf, read_rf_p1, 
         read_rf_p2, rtype_itypen, compute_sext, jump_sext : out std_logic;  
         alu_op_type : out std_logic_vector (3 downto 0);  sel_val_a, sel_val_b
         , signed_notsigned, alu_cin : out std_logic;  evaluate_branch : out 
         std_logic_vector (1 downto 0);  alu_overflow, zero_mul_detect, 
         mul_exeception : in std_logic;  dram_enable_cu, dram_r_nw_cu : out 
         std_logic;  dram_ready_cu : in std_logic;  update_pc_branch, write_rf,
         select_wb : out std_logic);

end control_unit_PC_SIZE32_RF_REGS32_IR_SIZE32_CW_SIZE22;

architecture SYN_behavioural of 
   control_unit_PC_SIZE32_RF_REGS32_IR_SIZE32_CW_SIZE22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component reg_nbit_n22_1
      port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0); 
            Q : out std_logic_vector (21 downto 0));
   end component;
   
   component reg_nbit_n22_2
      port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0); 
            Q : out std_logic_vector (21 downto 0));
   end component;
   
   component reg_nbit_n22_0
      port( clk, reset : in std_logic;  d : in std_logic_vector (21 downto 0); 
            Q : out std_logic_vector (21 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal stall_pip_port, enable_rf_port, read_rf_p2_port, rtype_itypen_port, 
      compute_sext_port, jump_sext_port, next_val_counter_mul_3_port, 
      next_val_counter_mul_2_port, next_val_counter_mul_1_port, 
      next_val_counter_mul_0_port, next_stall, cmd_word_17, cmd_word_8_port, 
      cmd_word_7_port, cmd_word_6_port, cmd_word_4_port, cmd_word_3_port, 
      cmd_word_2_port, cmd_word_1_port, cmd_alu_op_type_3_port, 
      cmd_alu_op_type_2_port, cmd_alu_op_type_1_port, cmd_alu_op_type_0_port, 
      N264, N265, N266, N267, N273, N274, N275, N276, N277, N278, N279, 
      cw1_21_port, cw1_20_port, cw1_19_port, cw1_18_port, cw1_17_port, 
      cw1_16_port, cw1_15_port, cw1_14_port, cw1_13_port, cw1_12_port, 
      cw1_11_port, cw1_10_port, cw1_9_port, cw1_8_port, cw1_7_port, cw1_6_port,
      cw1_5_port, cw1_4_port, cw1_3_port, cw1_2_port, cw1_1_port, cw1_0_port, 
      cw2_21_port, cw2_20_port, cw2_19_port, cw2_18_port, cw2_17_port, 
      cw2_16_port, cw2_15_port, cw2_14_port, cw2_13_port, cw2_12_port, 
      cw2_11_port, cw2_10_port, cw2_9_port, cw2_8_port, cw2_7_port, cw2_6_port,
      cw2_5_port, cw2_4_port, cw2_3_port, cw2_2_port, cw2_1_port, cw2_0_port, 
      cw3_21_port, cw3_20_port, cw3_19_port, cw3_18_port, cw3_17_port, 
      cw3_16_port, cw3_15_port, cw3_14_port, cw3_13_port, cw3_12_port, 
      cw3_11_port, cw3_10_port, cw3_9_port, cw3_8_port, cw3_7_port, cw3_6_port,
      cw3_5_port, cw3_4_port, cw3_3_port, cw3_2_port, cw3_1_port, cw3_0_port, 
      cw1_i_21_port, cw1_i_20_port, cw1_i_19_port, cw1_i_18_port, cw1_i_17_port
      , cw1_i_16_port, cw1_i_15_port, cw1_i_14_port, cw1_i_13_port, 
      cw1_i_12_port, cw1_i_11_port, cw1_i_9_port, cw1_i_8_port, cw1_i_7_port, 
      cw1_i_4_port, cw1_i_3_port, cw1_i_2_port, cw1_i_1_port, cw1_i_0_port, 
      cw2_i_21_port, cw2_i_20_port, cw2_i_19_port, cw2_i_18_port, cw2_i_17_port
      , cw2_i_16_port, cw2_i_15_port, cw2_i_14_port, cw2_i_13_port, 
      cw2_i_12_port, cw2_i_11_port, cw2_i_10_port, cw2_i_9_port, cw2_i_8_port, 
      cw2_i_7_port, cw2_i_4_port, cw2_i_3_port, cw2_i_2_port, cw2_i_1_port, 
      cw2_i_0_port, n23, n25, n26, n145, n209, n210, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n24, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n131, n132, n133, n134, n135, 
      n_5538, n_5539, n_5540 : std_logic;

begin
   stall_pip <= stall_pip_port;
   enable_rf <= enable_rf_port;
   read_rf_p1 <= enable_rf_port;
   read_rf_p2 <= read_rf_p2_port;
   rtype_itypen <= rtype_itypen_port;
   compute_sext <= compute_sext_port;
   jump_sext <= jump_sext_port;
   
   curr_state_reg_0_inst : DFFS_X1 port map( D => n210, CK => n6, SN => rst, Q 
                           => n2, QN => n23);
   curr_state_reg_1_inst : DFFR_X1 port map( D => n209, CK => n6, RN => rst, Q 
                           => n_5538, QN => n123);
   next_stall_reg : DLH_X1 port map( G => N279, D => n145, Q => next_stall);
   next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => N274, D => N273, Q 
                           => next_val_counter_mul_0_port);
   counter_mul_reg_0_inst : DFFR_X1 port map( D => next_val_counter_mul_0_port,
                           CK => n6, RN => rst, Q => n_5539, QN => n125);
   next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => N274, D => N277, Q 
                           => next_val_counter_mul_3_port);
   counter_mul_reg_3_inst : DFFR_X1 port map( D => next_val_counter_mul_3_port,
                           CK => n6, RN => rst, Q => n_5540, QN => n124);
   next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => N274, D => N276, Q 
                           => next_val_counter_mul_2_port);
   counter_mul_reg_2_inst : DFFR_X1 port map( D => next_val_counter_mul_2_port,
                           CK => n6, RN => rst, Q => n1, QN => n25);
   next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => N274, D => N275, Q 
                           => next_val_counter_mul_1_port);
   counter_mul_reg_1_inst : DFFR_X1 port map( D => next_val_counter_mul_1_port,
                           CK => n6, RN => rst, Q => n3, QN => n26);
   cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => N278, D => N267, Q => 
                           cmd_alu_op_type_3_port);
   cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => N278, D => N266, Q => 
                           cmd_alu_op_type_2_port);
   cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => N278, D => N265, Q => 
                           cmd_alu_op_type_1_port);
   cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => N278, D => N264, Q => 
                           cmd_alu_op_type_0_port);
   e_reg : reg_nbit_n22_0 port map( clk => n6, reset => n135, d(21) => 
                           cmd_word_17, d(20) => enable_rf_port, d(19) => 
                           enable_rf_port, d(18) => read_rf_p2_port, d(17) => 
                           rtype_itypen_port, d(16) => compute_sext_port, d(15)
                           => jump_sext_port, d(14) => n134, d(13) => 
                           compute_sext_port, d(12) => cmd_word_8_port, d(11) 
                           => cmd_word_7_port, d(10) => cmd_word_6_port, d(9) 
                           => n133, d(8) => cmd_word_4_port, d(7) => 
                           cmd_word_3_port, d(6) => cmd_word_2_port, d(5) => 
                           cmd_word_1_port, d(4) => n134, d(3) => 
                           cmd_alu_op_type_3_port, d(2) => 
                           cmd_alu_op_type_2_port, d(1) => 
                           cmd_alu_op_type_1_port, d(0) => 
                           cmd_alu_op_type_0_port, Q(21) => cw1_21_port, Q(20) 
                           => cw1_20_port, Q(19) => cw1_19_port, Q(18) => 
                           cw1_18_port, Q(17) => cw1_17_port, Q(16) => 
                           cw1_16_port, Q(15) => cw1_15_port, Q(14) => 
                           cw1_14_port, Q(13) => cw1_13_port, Q(12) => 
                           cw1_12_port, Q(11) => cw1_11_port, Q(10) => 
                           cw1_10_port, Q(9) => cw1_9_port, Q(8) => cw1_8_port,
                           Q(7) => cw1_7_port, Q(6) => cw1_6_port, Q(5) => 
                           cw1_5_port, Q(4) => cw1_4_port, Q(3) => cw1_3_port, 
                           Q(2) => cw1_2_port, Q(1) => cw1_1_port, Q(0) => 
                           cw1_0_port);
   m_reg : reg_nbit_n22_2 port map( clk => n6, reset => n135, d(21) => 
                           cw1_i_21_port, d(20) => cw1_i_20_port, d(19) => 
                           cw1_i_19_port, d(18) => cw1_i_18_port, d(17) => 
                           cw1_i_17_port, d(16) => cw1_i_16_port, d(15) => 
                           cw1_i_15_port, d(14) => cw1_i_14_port, d(13) => 
                           cw1_i_13_port, d(12) => cw1_i_12_port, d(11) => 
                           cw1_i_11_port, d(10) => n128, d(9) => cw1_i_9_port, 
                           d(8) => cw1_i_8_port, d(7) => cw1_i_7_port, d(6) => 
                           n127, d(5) => n126, d(4) => cw1_i_4_port, d(3) => 
                           cw1_i_3_port, d(2) => cw1_i_2_port, d(1) => 
                           cw1_i_1_port, d(0) => cw1_i_0_port, Q(21) => 
                           cw2_21_port, Q(20) => cw2_20_port, Q(19) => 
                           cw2_19_port, Q(18) => cw2_18_port, Q(17) => 
                           cw2_17_port, Q(16) => cw2_16_port, Q(15) => 
                           cw2_15_port, Q(14) => cw2_14_port, Q(13) => 
                           cw2_13_port, Q(12) => cw2_12_port, Q(11) => 
                           cw2_11_port, Q(10) => cw2_10_port, Q(9) => 
                           cw2_9_port, Q(8) => cw2_8_port, Q(7) => cw2_7_port, 
                           Q(6) => cw2_6_port, Q(5) => cw2_5_port, Q(4) => 
                           cw2_4_port, Q(3) => cw2_3_port, Q(2) => cw2_2_port, 
                           Q(1) => cw2_1_port, Q(0) => cw2_0_port);
   wb_reg : reg_nbit_n22_1 port map( clk => n6, reset => n135, d(21) => 
                           cw2_i_21_port, d(20) => cw2_i_20_port, d(19) => 
                           cw2_i_19_port, d(18) => cw2_i_18_port, d(17) => 
                           cw2_i_17_port, d(16) => cw2_i_16_port, d(15) => 
                           cw2_i_15_port, d(14) => cw2_i_14_port, d(13) => 
                           cw2_i_13_port, d(12) => cw2_i_12_port, d(11) => 
                           cw2_i_11_port, d(10) => cw2_i_10_port, d(9) => 
                           cw2_i_9_port, d(8) => cw2_i_8_port, d(7) => 
                           cw2_i_7_port, d(6) => n132, d(5) => n131, d(4) => 
                           cw2_i_4_port, d(3) => cw2_i_3_port, d(2) => 
                           cw2_i_2_port, d(1) => cw2_i_1_port, d(0) => 
                           cw2_i_0_port, Q(21) => cw3_21_port, Q(20) => 
                           cw3_20_port, Q(19) => cw3_19_port, Q(18) => 
                           cw3_18_port, Q(17) => cw3_17_port, Q(16) => 
                           cw3_16_port, Q(15) => cw3_15_port, Q(14) => 
                           cw3_14_port, Q(13) => cw3_13_port, Q(12) => 
                           cw3_12_port, Q(11) => cw3_11_port, Q(10) => 
                           cw3_10_port, Q(9) => cw3_9_port, Q(8) => cw3_8_port,
                           Q(7) => cw3_7_port, Q(6) => cw3_6_port, Q(5) => 
                           cw3_5_port, Q(4) => cw3_4_port, Q(3) => cw3_3_port, 
                           Q(2) => cw3_2_port, Q(1) => cw3_1_port, Q(0) => 
                           cw3_0_port);
   stall_reg : DFFR_X2 port map( D => next_stall, CK => n6, RN => rst, Q => 
                           stall_pip_port, QN => n4);
   U3 : INV_X4 port map( A => rst, ZN => n135);
   U4 : MUX2_X2 port map( A => cw1_14_port, B => n134, S => stall_pip_port, Z 
                           => sel_val_a);
   U5 : MUX2_X2 port map( A => cw1_13_port, B => compute_sext_port, S => 
                           stall_pip_port, Z => sel_val_b);
   U6 : INV_X2 port map( A => n17, ZN => compute_sext_port);
   U7 : OAI21_X4 port map( B1 => n7, B2 => n8, A => n10, ZN => select_wb);
   U8 : INV_X4 port map( A => n4, ZN => n5);
   U9 : BUF_X1 port map( A => clk, Z => n6);
   U10 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => write_rf);
   U11 : INV_X1 port map( A => cw3_5_port, ZN => n9);
   U12 : MUX2_X1 port map( A => cw2_4_port, B => n134, S => stall_pip_port, Z 
                           => update_pc_branch);
   U13 : MUX2_X1 port map( A => cw1_9_port, B => n133, S => stall_pip_port, Z 
                           => signed_notsigned);
   U14 : INV_X1 port map( A => cw3_6_port, ZN => n10);
   U15 : INV_X1 port map( A => n11, ZN => rtype_itypen_port);
   U16 : OR4_X1 port map( A1 => n12, A2 => cmd_word_3_port, A3 => 
                           cmd_word_7_port, A4 => read_rf_p2_port, ZN => 
                           enable_rf_port);
   U17 : OAI21_X1 port map( B1 => n13, B2 => n14, A => n11, ZN => 
                           read_rf_p2_port);
   U18 : AOI21_X1 port map( B1 => n15, B2 => n16, A => n13, ZN => n12);
   U19 : MUX2_X1 port map( A => cw1_5_port, B => cw2_5_port, S => 
                           stall_pip_port, Z => n126);
   U20 : MUX2_X1 port map( A => cw1_6_port, B => cw2_6_port, S => 
                           stall_pip_port, Z => n127);
   U21 : MUX2_X1 port map( A => cw1_10_port, B => cw2_10_port, S => 
                           stall_pip_port, Z => n128);
   U22 : MUX2_X1 port map( A => cw1_10_port, B => cmd_word_6_port, S => 
                           stall_pip_port, Z => evaluate_branch(0));
   U23 : MUX2_X1 port map( A => cw2_5_port, B => cw3_5_port, S => 
                           stall_pip_port, Z => n131);
   U24 : MUX2_X1 port map( A => cw2_6_port, B => cw3_6_port, S => 
                           stall_pip_port, Z => n132);
   U25 : NAND2_X1 port map( A1 => n11, A2 => n17, ZN => n133);
   U26 : OAI21_X1 port map( B1 => n18, B2 => n19, A => n20, ZN => n11);
   U27 : NOR2_X1 port map( A1 => n123, A2 => n23, ZN => n210);
   U28 : OR3_X1 port map( A1 => cmd_word_4_port, A2 => n134, A3 => n21, ZN => 
                           n209);
   U29 : INV_X1 port map( A => n22, ZN => n21);
   U30 : AOI22_X1 port map( A1 => n24, A2 => n27, B1 => n123, B2 => n2, ZN => 
                           n22);
   U31 : OAI21_X1 port map( B1 => n16, B2 => n28, A => n29, ZN => n27);
   U32 : MUX2_X1 port map( A => n30, B => n31, S => n32, Z => n29);
   U33 : NOR4_X1 port map( A1 => n33, A2 => curr_instruction_to_cu(13), A3 => 
                           curr_instruction_to_cu(15), A4 => 
                           curr_instruction_to_cu(14), ZN => n31);
   U34 : OR2_X1 port map( A1 => curr_instruction_to_cu(12), A2 => 
                           curr_instruction_to_cu(11), ZN => n33);
   U35 : NOR4_X1 port map( A1 => n34, A2 => curr_instruction_to_cu(18), A3 => 
                           curr_instruction_to_cu(20), A4 => 
                           curr_instruction_to_cu(19), ZN => n28);
   U36 : OR2_X1 port map( A1 => curr_instruction_to_cu(17), A2 => 
                           curr_instruction_to_cu(16), ZN => n34);
   U37 : NOR2_X1 port map( A1 => n13, A2 => n35, ZN => n134);
   U38 : NOR2_X1 port map( A1 => n5, A2 => n36, ZN => iram_enable_cu);
   U39 : INV_X1 port map( A => cmd_word_17, ZN => n36);
   U40 : MUX2_X1 port map( A => cw1_11_port, B => cmd_word_7_port, S => n5, Z 
                           => evaluate_branch(1));
   U41 : MUX2_X1 port map( A => cw2_7_port, B => cmd_word_3_port, S => n5, Z =>
                           dram_r_nw_cu);
   U42 : MUX2_X1 port map( A => cw2_8_port, B => cmd_word_4_port, S => n5, Z =>
                           dram_enable_cu);
   U43 : MUX2_X1 port map( A => cw2_9_port, B => cw3_9_port, S => n5, Z => 
                           cw2_i_9_port);
   U44 : MUX2_X1 port map( A => cw2_8_port, B => cw3_8_port, S => n5, Z => 
                           cw2_i_8_port);
   U45 : MUX2_X1 port map( A => cw2_7_port, B => cw3_7_port, S => n5, Z => 
                           cw2_i_7_port);
   U46 : MUX2_X1 port map( A => cw2_4_port, B => cw3_4_port, S => n5, Z => 
                           cw2_i_4_port);
   U47 : MUX2_X1 port map( A => cw2_3_port, B => cw3_3_port, S => n5, Z => 
                           cw2_i_3_port);
   U48 : MUX2_X1 port map( A => cw2_2_port, B => cw3_2_port, S => n5, Z => 
                           cw2_i_2_port);
   U49 : MUX2_X1 port map( A => cw2_21_port, B => cw3_21_port, S => n5, Z => 
                           cw2_i_21_port);
   U50 : MUX2_X1 port map( A => cw2_20_port, B => cw3_20_port, S => n5, Z => 
                           cw2_i_20_port);
   U51 : MUX2_X1 port map( A => cw2_1_port, B => cw3_1_port, S => n5, Z => 
                           cw2_i_1_port);
   U52 : MUX2_X1 port map( A => cw2_19_port, B => cw3_19_port, S => n5, Z => 
                           cw2_i_19_port);
   U53 : MUX2_X1 port map( A => cw2_18_port, B => cw3_18_port, S => n5, Z => 
                           cw2_i_18_port);
   U54 : MUX2_X1 port map( A => cw2_17_port, B => cw3_17_port, S => n5, Z => 
                           cw2_i_17_port);
   U55 : MUX2_X1 port map( A => cw2_16_port, B => cw3_16_port, S => n5, Z => 
                           cw2_i_16_port);
   U56 : MUX2_X1 port map( A => cw2_15_port, B => cw3_15_port, S => n5, Z => 
                           cw2_i_15_port);
   U57 : MUX2_X1 port map( A => cw2_14_port, B => cw3_14_port, S => n5, Z => 
                           cw2_i_14_port);
   U58 : MUX2_X1 port map( A => cw2_13_port, B => cw3_13_port, S => n5, Z => 
                           cw2_i_13_port);
   U59 : MUX2_X1 port map( A => cw2_12_port, B => cw3_12_port, S => n5, Z => 
                           cw2_i_12_port);
   U60 : MUX2_X1 port map( A => cw2_11_port, B => cw3_11_port, S => n5, Z => 
                           cw2_i_11_port);
   U61 : MUX2_X1 port map( A => cw2_10_port, B => cw3_10_port, S => n5, Z => 
                           cw2_i_10_port);
   U62 : MUX2_X1 port map( A => cw2_0_port, B => cw3_0_port, S => n5, Z => 
                           cw2_i_0_port);
   U63 : MUX2_X1 port map( A => cw1_9_port, B => cw2_9_port, S => n5, Z => 
                           cw1_i_9_port);
   U64 : MUX2_X1 port map( A => cw1_8_port, B => cw2_8_port, S => n5, Z => 
                           cw1_i_8_port);
   U65 : MUX2_X1 port map( A => cw1_7_port, B => cw2_7_port, S => n5, Z => 
                           cw1_i_7_port);
   U66 : MUX2_X1 port map( A => cw1_4_port, B => cw2_4_port, S => n5, Z => 
                           cw1_i_4_port);
   U67 : MUX2_X1 port map( A => cw1_3_port, B => cw2_3_port, S => n5, Z => 
                           cw1_i_3_port);
   U68 : MUX2_X1 port map( A => cw1_2_port, B => cw2_2_port, S => n5, Z => 
                           cw1_i_2_port);
   U69 : MUX2_X1 port map( A => cw1_21_port, B => cw2_21_port, S => n5, Z => 
                           cw1_i_21_port);
   U70 : MUX2_X1 port map( A => cw1_20_port, B => cw2_20_port, S => n5, Z => 
                           cw1_i_20_port);
   U71 : MUX2_X1 port map( A => cw1_1_port, B => cw2_1_port, S => n5, Z => 
                           cw1_i_1_port);
   U72 : MUX2_X1 port map( A => cw1_19_port, B => cw2_19_port, S => n5, Z => 
                           cw1_i_19_port);
   U73 : MUX2_X1 port map( A => cw1_18_port, B => cw2_18_port, S => n5, Z => 
                           cw1_i_18_port);
   U74 : MUX2_X1 port map( A => cw1_17_port, B => cw2_17_port, S => n5, Z => 
                           cw1_i_17_port);
   U75 : MUX2_X1 port map( A => cw1_16_port, B => cw2_16_port, S => n5, Z => 
                           cw1_i_16_port);
   U76 : MUX2_X1 port map( A => cw1_15_port, B => cw2_15_port, S => n5, Z => 
                           cw1_i_15_port);
   U77 : MUX2_X1 port map( A => cw1_14_port, B => cw2_14_port, S => n5, Z => 
                           cw1_i_14_port);
   U78 : MUX2_X1 port map( A => cw1_13_port, B => cw2_13_port, S => n5, Z => 
                           cw1_i_13_port);
   U79 : MUX2_X1 port map( A => cw1_12_port, B => cw2_12_port, S => n5, Z => 
                           cw1_i_12_port);
   U80 : MUX2_X1 port map( A => cw1_11_port, B => cw2_11_port, S => n5, Z => 
                           cw1_i_11_port);
   U81 : MUX2_X1 port map( A => cw1_0_port, B => cw2_0_port, S => n5, Z => 
                           cw1_i_0_port);
   U82 : OAI211_X1 port map( C1 => n18, C2 => n37, A => n17, B => n38, ZN => 
                           cmd_word_17);
   U83 : AOI22_X1 port map( A1 => n24, A2 => n39, B1 => n123, B2 => n2, ZN => 
                           n38);
   U84 : OAI21_X1 port map( B1 => n40, B2 => n41, A => n42, ZN => n39);
   U85 : MUX2_X1 port map( A => n5, B => n43, S => n32, Z => n42);
   U86 : AND2_X1 port map( A1 => n145, A2 => n7, ZN => n18);
   U87 : INV_X1 port map( A => n44, ZN => n7);
   U88 : NOR2_X1 port map( A1 => n45, A2 => n13, ZN => cmd_word_7_port);
   U89 : OAI21_X1 port map( B1 => n13, B2 => n15, A => n46, ZN => 
                           cmd_word_6_port);
   U90 : INV_X1 port map( A => jump_sext_port, ZN => n46);
   U91 : NOR2_X1 port map( A1 => n13, A2 => n47, ZN => jump_sext_port);
   U92 : OAI21_X1 port map( B1 => n13, B2 => n14, A => n48, ZN => 
                           cmd_word_4_port);
   U93 : INV_X1 port map( A => n49, ZN => cmd_word_2_port);
   U94 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => cmd_word_1_port);
   U95 : OAI21_X1 port map( B1 => n50, B2 => n51, A => n24, ZN => n49);
   U96 : OAI21_X1 port map( B1 => n43, B2 => n52, A => n53, ZN => n51);
   U97 : INV_X1 port map( A => cmd_word_3_port, ZN => n48);
   U98 : NOR2_X1 port map( A1 => n54, A2 => n13, ZN => cmd_word_3_port);
   U99 : MUX2_X1 port map( A => cw1_3_port, B => cmd_alu_op_type_3_port, S => 
                           n5, Z => alu_op_type(3));
   U100 : MUX2_X1 port map( A => cw1_2_port, B => cmd_alu_op_type_2_port, S => 
                           n5, Z => alu_op_type(2));
   U101 : MUX2_X1 port map( A => cw1_1_port, B => cmd_alu_op_type_1_port, S => 
                           n5, Z => alu_op_type(1));
   U102 : MUX2_X1 port map( A => cw1_0_port, B => cmd_alu_op_type_0_port, S => 
                           n5, Z => alu_op_type(0));
   U103 : MUX2_X1 port map( A => cw1_12_port, B => cmd_word_8_port, S => n5, Z 
                           => alu_cin);
   U104 : OAI22_X1 port map( A1 => n13, A2 => n55, B1 => n37, B2 => n56, ZN => 
                           cmd_word_8_port);
   U105 : INV_X1 port map( A => n24, ZN => n13);
   U106 : AOI211_X1 port map( C1 => n5, C2 => n145, A => n8, B => n44, ZN => 
                           N279);
   U107 : AOI21_X1 port map( B1 => n25, B2 => n26, A => n124, ZN => n44);
   U108 : OR4_X1 port map( A1 => n3, A2 => n1, A3 => n125, A4 => n124, ZN => 
                           n145);
   U109 : NAND2_X1 port map( A1 => n17, A2 => n37, ZN => N278);
   U110 : NAND2_X1 port map( A1 => n24, A2 => n30, ZN => n17);
   U111 : NAND4_X1 port map( A1 => n35, A2 => n16, A3 => n14, A4 => n54, ZN => 
                           n30);
   U112 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n54);
   U113 : NAND2_X1 port map( A1 => n57, A2 => curr_instruction_to_cu(29), ZN =>
                           n14);
   U114 : AND4_X1 port map( A1 => curr_instruction_to_cu(31), A2 => 
                           curr_instruction_to_cu(27), A3 => 
                           curr_instruction_to_cu(26), A4 => n59, ZN => n57);
   U115 : INV_X1 port map( A => n50, ZN => n16);
   U116 : OAI211_X1 port map( C1 => n40, C2 => n60, A => n61, B => n62, ZN => 
                           n50);
   U117 : AOI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n62);
   U118 : INV_X1 port map( A => n66, ZN => n65);
   U119 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n41, ZN => n64);
   U120 : INV_X1 port map( A => n69, ZN => n68);
   U121 : INV_X1 port map( A => n70, ZN => n40);
   U122 : AND3_X1 port map( A1 => n15, A2 => n45, A3 => n47, ZN => n35);
   U123 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n47);
   U124 : INV_X1 port map( A => n53, ZN => n73);
   U125 : NAND3_X1 port map( A1 => curr_instruction_to_cu(26), A2 => n71, A3 =>
                           curr_instruction_to_cu(27), ZN => n53);
   U126 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n70, ZN => n45);
   U127 : NAND3_X1 port map( A1 => n63, A2 => n75, A3 => n74, ZN => n15);
   U128 : MUX2_X1 port map( A => n76, B => n77, S => n124, Z => N277);
   U129 : NOR3_X1 port map( A1 => n78, A2 => n26, A3 => n25, ZN => n77);
   U130 : OAI21_X1 port map( B1 => n1, B2 => n8, A => n79, ZN => n76);
   U131 : MUX2_X1 port map( A => n80, B => n81, S => n25, Z => N276);
   U132 : NOR2_X1 port map( A1 => n26, A2 => n78, ZN => n81);
   U133 : INV_X1 port map( A => n82, ZN => n78);
   U134 : INV_X1 port map( A => n79, ZN => n80);
   U135 : AOI21_X1 port map( B1 => n26, B2 => n83, A => N273, ZN => n79);
   U136 : MUX2_X1 port map( A => N273, B => n82, S => n26, Z => N275);
   U137 : NOR2_X1 port map( A1 => n8, A2 => n125, ZN => n82);
   U138 : NAND2_X1 port map( A1 => n5, A2 => n8, ZN => N274);
   U139 : AND2_X1 port map( A1 => n125, A2 => n83, ZN => N273);
   U140 : INV_X1 port map( A => n8, ZN => n83);
   U141 : NAND2_X1 port map( A1 => n20, A2 => n43, ZN => n8);
   U142 : INV_X1 port map( A => n37, ZN => n20);
   U143 : NAND2_X1 port map( A1 => n32, A2 => n24, ZN => n37);
   U144 : NOR2_X1 port map( A1 => n2, A2 => n123, ZN => n24);
   U145 : NAND3_X1 port map( A1 => n66, A2 => n84, A3 => n85, ZN => N267);
   U146 : OR3_X1 port map( A1 => n52, A2 => n86, A3 => n87, ZN => n85);
   U147 : NAND3_X1 port map( A1 => n69, A2 => n70, A3 => 
                           curr_instruction_to_cu(30), ZN => n66);
   U148 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n90, ZN => N266);
   U149 : NAND3_X1 port map( A1 => n32, A2 => n91, A3 => n92, ZN => n89);
   U150 : INV_X1 port map( A => n93, ZN => n92);
   U151 : XOR2_X1 port map( A => curr_instruction_to_cu(1), B => 
                           curr_instruction_to_cu(0), Z => n91);
   U152 : OAI21_X1 port map( B1 => n70, B2 => n72, A => n94, ZN => n88);
   U153 : NAND4_X1 port map( A1 => n90, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           N265);
   U154 : NAND4_X1 port map( A1 => curr_instruction_to_cu(30), A2 => n69, A3 =>
                           n70, A4 => n98, ZN => n97);
   U155 : NOR2_X1 port map( A1 => n99, A2 => curr_instruction_to_cu(27), ZN => 
                           n70);
   U156 : OAI21_X1 port map( B1 => n43, B2 => n100, A => n32, ZN => n96);
   U157 : MUX2_X1 port map( A => n101, B => n102, S => 
                           curr_instruction_to_cu(0), Z => n100);
   U158 : NOR2_X1 port map( A1 => curr_instruction_to_cu(2), A2 => n87, ZN => 
                           n102);
   U159 : NOR2_X1 port map( A1 => curr_instruction_to_cu(1), A2 => n93, ZN => 
                           n101);
   U160 : INV_X1 port map( A => n19, ZN => n43);
   U161 : NAND4_X1 port map( A1 => curr_instruction_to_cu(1), A2 => 
                           curr_instruction_to_cu(0), A3 => 
                           curr_instruction_to_cu(2), A4 => n103, ZN => n19);
   U162 : AND3_X1 port map( A1 => curr_instruction_to_cu(5), A2 => 
                           curr_instruction_to_cu(3), A3 => 
                           curr_instruction_to_cu(4), ZN => n103);
   U163 : NAND2_X1 port map( A1 => n94, A2 => n63, ZN => n95);
   U164 : INV_X1 port map( A => n60, ZN => n94);
   U165 : INV_X1 port map( A => n104, ZN => n90);
   U166 : OAI21_X1 port map( B1 => n105, B2 => n41, A => n106, ZN => n104);
   U167 : NAND4_X1 port map( A1 => n32, A2 => n107, A3 => 
                           curr_instruction_to_cu(2), A4 => n108, ZN => n106);
   U168 : NOR3_X1 port map( A1 => curr_instruction_to_cu(3), A2 => 
                           curr_instruction_to_cu(5), A3 => 
                           curr_instruction_to_cu(4), ZN => n108);
   U169 : INV_X1 port map( A => n52, ZN => n32);
   U170 : OAI21_X1 port map( B1 => n109, B2 => n52, A => n61, ZN => N264);
   U171 : AND3_X1 port map( A1 => n84, A2 => n55, A3 => n110, ZN => n61);
   U172 : INV_X1 port map( A => n111, ZN => n110);
   U173 : OAI22_X1 port map( A1 => n60, A2 => n105, B1 => n41, B2 => n112, ZN 
                           => n111);
   U174 : NAND2_X1 port map( A1 => curr_instruction_to_cu(30), A2 => n74, ZN =>
                           n41);
   U175 : NOR3_X1 port map( A1 => curr_instruction_to_cu(29), A2 => 
                           curr_instruction_to_cu(31), A3 => n98, ZN => n74);
   U176 : NOR2_X1 port map( A1 => n63, A2 => n72, ZN => n105);
   U177 : NAND3_X1 port map( A1 => curr_instruction_to_cu(28), A2 => n75, A3 =>
                           n69, ZN => n60);
   U178 : NAND3_X1 port map( A1 => n72, A2 => n59, A3 => n69, ZN => n55);
   U179 : INV_X1 port map( A => n67, ZN => n59);
   U180 : INV_X1 port map( A => n112, ZN => n72);
   U181 : NAND2_X1 port map( A1 => curr_instruction_to_cu(27), A2 => n99, ZN =>
                           n112);
   U182 : INV_X1 port map( A => curr_instruction_to_cu(26), ZN => n99);
   U183 : NAND4_X1 port map( A1 => curr_instruction_to_cu(30), A2 => n69, A3 =>
                           curr_instruction_to_cu(28), A4 => n63, ZN => n84);
   U184 : NOR2_X1 port map( A1 => n58, A2 => curr_instruction_to_cu(31), ZN => 
                           n69);
   U185 : INV_X1 port map( A => curr_instruction_to_cu(29), ZN => n58);
   U186 : NAND2_X1 port map( A1 => n71, A2 => n63, ZN => n52);
   U187 : NOR2_X1 port map( A1 => curr_instruction_to_cu(26), A2 => 
                           curr_instruction_to_cu(27), ZN => n63);
   U188 : NOR3_X1 port map( A1 => curr_instruction_to_cu(29), A2 => 
                           curr_instruction_to_cu(31), A3 => n67, ZN => n71);
   U189 : NAND2_X1 port map( A1 => n98, A2 => n75, ZN => n67);
   U190 : INV_X1 port map( A => curr_instruction_to_cu(30), ZN => n75);
   U191 : INV_X1 port map( A => curr_instruction_to_cu(28), ZN => n98);
   U192 : AOI21_X1 port map( B1 => n113, B2 => n107, A => n114, ZN => n109);
   U193 : INV_X1 port map( A => n56, ZN => n114);
   U194 : NAND3_X1 port map( A1 => n115, A2 => curr_instruction_to_cu(1), A3 =>
                           n86, ZN => n56);
   U195 : NOR2_X1 port map( A1 => curr_instruction_to_cu(2), A2 => 
                           curr_instruction_to_cu(0), ZN => n86);
   U196 : INV_X1 port map( A => curr_instruction_to_cu(0), ZN => n107);
   U197 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n93, ZN => n113);
   U198 : NAND2_X1 port map( A1 => n115, A2 => curr_instruction_to_cu(2), ZN =>
                           n93);
   U199 : NOR3_X1 port map( A1 => curr_instruction_to_cu(3), A2 => 
                           curr_instruction_to_cu(4), A3 => n118, ZN => n115);
   U200 : INV_X1 port map( A => curr_instruction_to_cu(5), ZN => n118);
   U201 : INV_X1 port map( A => curr_instruction_to_cu(2), ZN => n117);
   U202 : NOR2_X1 port map( A1 => n119, A2 => n120, ZN => n116);
   U203 : INV_X1 port map( A => n87, ZN => n120);
   U204 : NAND4_X1 port map( A1 => curr_instruction_to_cu(5), A2 => 
                           curr_instruction_to_cu(3), A3 => n121, A4 => n122, 
                           ZN => n87);
   U205 : INV_X1 port map( A => curr_instruction_to_cu(4), ZN => n122);
   U206 : NOR3_X1 port map( A1 => n121, A2 => curr_instruction_to_cu(4), A3 => 
                           curr_instruction_to_cu(3), ZN => n119);
   U207 : INV_X1 port map( A => curr_instruction_to_cu(1), ZN => n121);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component DATAPATH_N32_RF_REGS32_IR_SIZE32_PC_SIZE32
      port( clk, rst : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
            downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic
            ;  IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : 
            out std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE
            : out std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
            std_logic_vector (31 downto 0);  iram_enable_cu : in std_logic;  
            iram_ready_cu : out std_logic;  stall : in std_logic;  
            curr_instruction_to_cu : out std_logic_vector (31 downto 0);  
            enable_rf, read_rf_p1, read_rf_p2, write_rf, rtype_itypen, 
            compute_sext, jump_sext : in std_logic;  alu_op_type : in 
            std_logic_vector (3 downto 0);  sel_val_a, sel_val_b, 
            signed_notsigned : in std_logic;  evaluate_branch : in 
            std_logic_vector (1 downto 0);  alu_cin : in std_logic;  
            alu_overflow, zero_mul_detect, mul_exeception : out std_logic;  
            dram_enable_cu, dram_r_nw_cu : in std_logic;  dram_ready_cu : out 
            std_logic;  update_pc_branch, select_wb : in std_logic);
   end component;
   
   component control_unit_PC_SIZE32_RF_REGS32_IR_SIZE32_CW_SIZE22
      port( clk, rst : in std_logic;  iram_enable_cu : out std_logic;  
            iram_ready_cu : in std_logic;  curr_instruction_to_cu : in 
            std_logic_vector (31 downto 0);  stall_pip, enable_rf, read_rf_p1, 
            read_rf_p2, rtype_itypen, compute_sext, jump_sext : out std_logic; 
            alu_op_type : out std_logic_vector (3 downto 0);  sel_val_a, 
            sel_val_b, signed_notsigned, alu_cin : out std_logic;  
            evaluate_branch : out std_logic_vector (1 downto 0);  alu_overflow,
            zero_mul_detect, mul_exeception : in std_logic;  dram_enable_cu, 
            dram_r_nw_cu : out std_logic;  dram_ready_cu : in std_logic;  
            update_pc_branch, write_rf, select_wb : out std_logic);
   end component;
   
   signal DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      iram_enable_cu_i, iram_ready_cu_i, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_29_port, 
      curr_instruction_to_cu_i_28_port, curr_instruction_to_cu_i_27_port, 
      curr_instruction_to_cu_i_26_port, curr_instruction_to_cu_i_25_port, 
      curr_instruction_to_cu_i_24_port, curr_instruction_to_cu_i_23_port, 
      curr_instruction_to_cu_i_22_port, curr_instruction_to_cu_i_21_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_10_port, curr_instruction_to_cu_i_9_port, 
      curr_instruction_to_cu_i_8_port, curr_instruction_to_cu_i_7_port, 
      curr_instruction_to_cu_i_6_port, curr_instruction_to_cu_i_5_port, 
      curr_instruction_to_cu_i_4_port, curr_instruction_to_cu_i_3_port, 
      curr_instruction_to_cu_i_2_port, curr_instruction_to_cu_i_1_port, 
      curr_instruction_to_cu_i_0_port, stall_i, enable_rf_i, read_rf_p1_i, 
      read_rf_p2_i, rtype_itypen_i, compute_sext_i, jump_sext_i, 
      alu_op_type_i_3_port, alu_op_type_i_2_port, alu_op_type_i_1_port, 
      alu_op_type_i_0_port, sel_val_a_i_0_port, sel_val_b_i_0_port, 
      signed_notsigned_i, alu_cin_i, evaluate_branch_i_1_port, 
      evaluate_branch_i_0_port, alu_overflow_i, zero_mul_detect_i, 
      mul_exeception_i, dram_enable_cu_i, dram_r_nw_cu_i, dram_ready_cu_i, 
      update_pc_branch_i, write_rf_i, select_wb_i_0_port, DRAM_ADDRESS_0_port, 
      n_5541, n_5542 : std_logic;

begin
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_0_port, DRAM_ADDRESS_0_port );
   
   cu_i : control_unit_PC_SIZE32_RF_REGS32_IR_SIZE32_CW_SIZE22 port map( clk =>
                           CLK, rst => RST, iram_enable_cu => iram_enable_cu_i,
                           iram_ready_cu => iram_ready_cu_i, 
                           curr_instruction_to_cu(31) => 
                           curr_instruction_to_cu_i_31_port, 
                           curr_instruction_to_cu(30) => 
                           curr_instruction_to_cu_i_30_port, 
                           curr_instruction_to_cu(29) => 
                           curr_instruction_to_cu_i_29_port, 
                           curr_instruction_to_cu(28) => 
                           curr_instruction_to_cu_i_28_port, 
                           curr_instruction_to_cu(27) => 
                           curr_instruction_to_cu_i_27_port, 
                           curr_instruction_to_cu(26) => 
                           curr_instruction_to_cu_i_26_port, 
                           curr_instruction_to_cu(25) => 
                           curr_instruction_to_cu_i_25_port, 
                           curr_instruction_to_cu(24) => 
                           curr_instruction_to_cu_i_24_port, 
                           curr_instruction_to_cu(23) => 
                           curr_instruction_to_cu_i_23_port, 
                           curr_instruction_to_cu(22) => 
                           curr_instruction_to_cu_i_22_port, 
                           curr_instruction_to_cu(21) => 
                           curr_instruction_to_cu_i_21_port, 
                           curr_instruction_to_cu(20) => 
                           curr_instruction_to_cu_i_20_port, 
                           curr_instruction_to_cu(19) => 
                           curr_instruction_to_cu_i_19_port, 
                           curr_instruction_to_cu(18) => 
                           curr_instruction_to_cu_i_18_port, 
                           curr_instruction_to_cu(17) => 
                           curr_instruction_to_cu_i_17_port, 
                           curr_instruction_to_cu(16) => 
                           curr_instruction_to_cu_i_16_port, 
                           curr_instruction_to_cu(15) => 
                           curr_instruction_to_cu_i_15_port, 
                           curr_instruction_to_cu(14) => 
                           curr_instruction_to_cu_i_14_port, 
                           curr_instruction_to_cu(13) => 
                           curr_instruction_to_cu_i_13_port, 
                           curr_instruction_to_cu(12) => 
                           curr_instruction_to_cu_i_12_port, 
                           curr_instruction_to_cu(11) => 
                           curr_instruction_to_cu_i_11_port, 
                           curr_instruction_to_cu(10) => 
                           curr_instruction_to_cu_i_10_port, 
                           curr_instruction_to_cu(9) => 
                           curr_instruction_to_cu_i_9_port, 
                           curr_instruction_to_cu(8) => 
                           curr_instruction_to_cu_i_8_port, 
                           curr_instruction_to_cu(7) => 
                           curr_instruction_to_cu_i_7_port, 
                           curr_instruction_to_cu(6) => 
                           curr_instruction_to_cu_i_6_port, 
                           curr_instruction_to_cu(5) => 
                           curr_instruction_to_cu_i_5_port, 
                           curr_instruction_to_cu(4) => 
                           curr_instruction_to_cu_i_4_port, 
                           curr_instruction_to_cu(3) => 
                           curr_instruction_to_cu_i_3_port, 
                           curr_instruction_to_cu(2) => 
                           curr_instruction_to_cu_i_2_port, 
                           curr_instruction_to_cu(1) => 
                           curr_instruction_to_cu_i_1_port, 
                           curr_instruction_to_cu(0) => 
                           curr_instruction_to_cu_i_0_port, stall_pip => 
                           stall_i, enable_rf => enable_rf_i, read_rf_p1 => 
                           read_rf_p1_i, read_rf_p2 => read_rf_p2_i, 
                           rtype_itypen => rtype_itypen_i, compute_sext => 
                           compute_sext_i, jump_sext => jump_sext_i, 
                           alu_op_type(3) => alu_op_type_i_3_port, 
                           alu_op_type(2) => alu_op_type_i_2_port, 
                           alu_op_type(1) => alu_op_type_i_1_port, 
                           alu_op_type(0) => alu_op_type_i_0_port, sel_val_a =>
                           sel_val_a_i_0_port, sel_val_b => sel_val_b_i_0_port,
                           signed_notsigned => signed_notsigned_i, alu_cin => 
                           alu_cin_i, evaluate_branch(1) => 
                           evaluate_branch_i_1_port, evaluate_branch(0) => 
                           evaluate_branch_i_0_port, alu_overflow => 
                           alu_overflow_i, zero_mul_detect => zero_mul_detect_i
                           , mul_exeception => mul_exeception_i, dram_enable_cu
                           => dram_enable_cu_i, dram_r_nw_cu => dram_r_nw_cu_i,
                           dram_ready_cu => dram_ready_cu_i, update_pc_branch 
                           => update_pc_branch_i, write_rf => write_rf_i, 
                           select_wb => select_wb_i_0_port);
   datapath_i : DATAPATH_N32_RF_REGS32_IR_SIZE32_PC_SIZE32 port map( clk => CLK
                           , rst => RST, IRAM_ADDRESS(31) => IRAM_ADDRESS(31), 
                           IRAM_ADDRESS(30) => IRAM_ADDRESS(30), 
                           IRAM_ADDRESS(29) => IRAM_ADDRESS(29), 
                           IRAM_ADDRESS(28) => IRAM_ADDRESS(28), 
                           IRAM_ADDRESS(27) => IRAM_ADDRESS(27), 
                           IRAM_ADDRESS(26) => IRAM_ADDRESS(26), 
                           IRAM_ADDRESS(25) => IRAM_ADDRESS(25), 
                           IRAM_ADDRESS(24) => IRAM_ADDRESS(24), 
                           IRAM_ADDRESS(23) => IRAM_ADDRESS(23), 
                           IRAM_ADDRESS(22) => IRAM_ADDRESS(22), 
                           IRAM_ADDRESS(21) => IRAM_ADDRESS(21), 
                           IRAM_ADDRESS(20) => IRAM_ADDRESS(20), 
                           IRAM_ADDRESS(19) => IRAM_ADDRESS(19), 
                           IRAM_ADDRESS(18) => IRAM_ADDRESS(18), 
                           IRAM_ADDRESS(17) => IRAM_ADDRESS(17), 
                           IRAM_ADDRESS(16) => IRAM_ADDRESS(16), 
                           IRAM_ADDRESS(15) => IRAM_ADDRESS(15), 
                           IRAM_ADDRESS(14) => IRAM_ADDRESS(14), 
                           IRAM_ADDRESS(13) => IRAM_ADDRESS(13), 
                           IRAM_ADDRESS(12) => IRAM_ADDRESS(12), 
                           IRAM_ADDRESS(11) => IRAM_ADDRESS(11), 
                           IRAM_ADDRESS(10) => IRAM_ADDRESS(10), 
                           IRAM_ADDRESS(9) => IRAM_ADDRESS(9), IRAM_ADDRESS(8) 
                           => IRAM_ADDRESS(8), IRAM_ADDRESS(7) => 
                           IRAM_ADDRESS(7), IRAM_ADDRESS(6) => IRAM_ADDRESS(6),
                           IRAM_ADDRESS(5) => IRAM_ADDRESS(5), IRAM_ADDRESS(4) 
                           => IRAM_ADDRESS(4), IRAM_ADDRESS(3) => 
                           IRAM_ADDRESS(3), IRAM_ADDRESS(2) => IRAM_ADDRESS(2),
                           IRAM_ADDRESS(1) => IRAM_ADDRESS(1), IRAM_ADDRESS(0) 
                           => IRAM_ADDRESS(0), IRAM_ENABLE => IRAM_ENABLE, 
                           IRAM_READY => IRAM_READY, IRAM_DATA(31) => 
                           IRAM_DATA(31), IRAM_DATA(30) => IRAM_DATA(30), 
                           IRAM_DATA(29) => IRAM_DATA(29), IRAM_DATA(28) => 
                           IRAM_DATA(28), IRAM_DATA(27) => IRAM_DATA(27), 
                           IRAM_DATA(26) => IRAM_DATA(26), IRAM_DATA(25) => 
                           IRAM_DATA(25), IRAM_DATA(24) => IRAM_DATA(24), 
                           IRAM_DATA(23) => IRAM_DATA(23), IRAM_DATA(22) => 
                           IRAM_DATA(22), IRAM_DATA(21) => IRAM_DATA(21), 
                           IRAM_DATA(20) => IRAM_DATA(20), IRAM_DATA(19) => 
                           IRAM_DATA(19), IRAM_DATA(18) => IRAM_DATA(18), 
                           IRAM_DATA(17) => IRAM_DATA(17), IRAM_DATA(16) => 
                           IRAM_DATA(16), IRAM_DATA(15) => IRAM_DATA(15), 
                           IRAM_DATA(14) => IRAM_DATA(14), IRAM_DATA(13) => 
                           IRAM_DATA(13), IRAM_DATA(12) => IRAM_DATA(12), 
                           IRAM_DATA(11) => IRAM_DATA(11), IRAM_DATA(10) => 
                           IRAM_DATA(10), IRAM_DATA(9) => IRAM_DATA(9), 
                           IRAM_DATA(8) => IRAM_DATA(8), IRAM_DATA(7) => 
                           IRAM_DATA(7), IRAM_DATA(6) => IRAM_DATA(6), 
                           IRAM_DATA(5) => IRAM_DATA(5), IRAM_DATA(4) => 
                           IRAM_DATA(4), IRAM_DATA(3) => IRAM_DATA(3), 
                           IRAM_DATA(2) => IRAM_DATA(2), IRAM_DATA(1) => 
                           IRAM_DATA(1), IRAM_DATA(0) => IRAM_DATA(0), 
                           DRAM_ADDRESS(31) => DRAM_ADDRESS_31_port, 
                           DRAM_ADDRESS(30) => DRAM_ADDRESS_30_port, 
                           DRAM_ADDRESS(29) => DRAM_ADDRESS_29_port, 
                           DRAM_ADDRESS(28) => DRAM_ADDRESS_28_port, 
                           DRAM_ADDRESS(27) => DRAM_ADDRESS_27_port, 
                           DRAM_ADDRESS(26) => DRAM_ADDRESS_26_port, 
                           DRAM_ADDRESS(25) => DRAM_ADDRESS_25_port, 
                           DRAM_ADDRESS(24) => DRAM_ADDRESS_24_port, 
                           DRAM_ADDRESS(23) => DRAM_ADDRESS_23_port, 
                           DRAM_ADDRESS(22) => DRAM_ADDRESS_22_port, 
                           DRAM_ADDRESS(21) => DRAM_ADDRESS_21_port, 
                           DRAM_ADDRESS(20) => DRAM_ADDRESS_20_port, 
                           DRAM_ADDRESS(19) => DRAM_ADDRESS_19_port, 
                           DRAM_ADDRESS(18) => DRAM_ADDRESS_18_port, 
                           DRAM_ADDRESS(17) => DRAM_ADDRESS_17_port, 
                           DRAM_ADDRESS(16) => DRAM_ADDRESS_16_port, 
                           DRAM_ADDRESS(15) => DRAM_ADDRESS_15_port, 
                           DRAM_ADDRESS(14) => DRAM_ADDRESS_14_port, 
                           DRAM_ADDRESS(13) => DRAM_ADDRESS_13_port, 
                           DRAM_ADDRESS(12) => DRAM_ADDRESS_12_port, 
                           DRAM_ADDRESS(11) => DRAM_ADDRESS_11_port, 
                           DRAM_ADDRESS(10) => DRAM_ADDRESS_10_port, 
                           DRAM_ADDRESS(9) => DRAM_ADDRESS_9_port, 
                           DRAM_ADDRESS(8) => DRAM_ADDRESS_8_port, 
                           DRAM_ADDRESS(7) => DRAM_ADDRESS_7_port, 
                           DRAM_ADDRESS(6) => DRAM_ADDRESS_6_port, 
                           DRAM_ADDRESS(5) => DRAM_ADDRESS_5_port, 
                           DRAM_ADDRESS(4) => DRAM_ADDRESS_4_port, 
                           DRAM_ADDRESS(3) => DRAM_ADDRESS_3_port, 
                           DRAM_ADDRESS(2) => DRAM_ADDRESS_2_port, 
                           DRAM_ADDRESS(1) => n_5541, DRAM_ADDRESS(0) => n_5542
                           , DRAM_ENABLE => DRAM_ENABLE, DRAM_READNOTWRITE => 
                           DRAM_READNOTWRITE, DRAM_READY => DRAM_READY, 
                           DRAM_DATA(31) => DRAM_DATA(31), DRAM_DATA(30) => 
                           DRAM_DATA(30), DRAM_DATA(29) => DRAM_DATA(29), 
                           DRAM_DATA(28) => DRAM_DATA(28), DRAM_DATA(27) => 
                           DRAM_DATA(27), DRAM_DATA(26) => DRAM_DATA(26), 
                           DRAM_DATA(25) => DRAM_DATA(25), DRAM_DATA(24) => 
                           DRAM_DATA(24), DRAM_DATA(23) => DRAM_DATA(23), 
                           DRAM_DATA(22) => DRAM_DATA(22), DRAM_DATA(21) => 
                           DRAM_DATA(21), DRAM_DATA(20) => DRAM_DATA(20), 
                           DRAM_DATA(19) => DRAM_DATA(19), DRAM_DATA(18) => 
                           DRAM_DATA(18), DRAM_DATA(17) => DRAM_DATA(17), 
                           DRAM_DATA(16) => DRAM_DATA(16), DRAM_DATA(15) => 
                           DRAM_DATA(15), DRAM_DATA(14) => DRAM_DATA(14), 
                           DRAM_DATA(13) => DRAM_DATA(13), DRAM_DATA(12) => 
                           DRAM_DATA(12), DRAM_DATA(11) => DRAM_DATA(11), 
                           DRAM_DATA(10) => DRAM_DATA(10), DRAM_DATA(9) => 
                           DRAM_DATA(9), DRAM_DATA(8) => DRAM_DATA(8), 
                           DRAM_DATA(7) => DRAM_DATA(7), DRAM_DATA(6) => 
                           DRAM_DATA(6), DRAM_DATA(5) => DRAM_DATA(5), 
                           DRAM_DATA(4) => DRAM_DATA(4), DRAM_DATA(3) => 
                           DRAM_DATA(3), DRAM_DATA(2) => DRAM_DATA(2), 
                           DRAM_DATA(1) => DRAM_DATA(1), DRAM_DATA(0) => 
                           DRAM_DATA(0), iram_enable_cu => iram_enable_cu_i, 
                           iram_ready_cu => iram_ready_cu_i, stall => stall_i, 
                           curr_instruction_to_cu(31) => 
                           curr_instruction_to_cu_i_31_port, 
                           curr_instruction_to_cu(30) => 
                           curr_instruction_to_cu_i_30_port, 
                           curr_instruction_to_cu(29) => 
                           curr_instruction_to_cu_i_29_port, 
                           curr_instruction_to_cu(28) => 
                           curr_instruction_to_cu_i_28_port, 
                           curr_instruction_to_cu(27) => 
                           curr_instruction_to_cu_i_27_port, 
                           curr_instruction_to_cu(26) => 
                           curr_instruction_to_cu_i_26_port, 
                           curr_instruction_to_cu(25) => 
                           curr_instruction_to_cu_i_25_port, 
                           curr_instruction_to_cu(24) => 
                           curr_instruction_to_cu_i_24_port, 
                           curr_instruction_to_cu(23) => 
                           curr_instruction_to_cu_i_23_port, 
                           curr_instruction_to_cu(22) => 
                           curr_instruction_to_cu_i_22_port, 
                           curr_instruction_to_cu(21) => 
                           curr_instruction_to_cu_i_21_port, 
                           curr_instruction_to_cu(20) => 
                           curr_instruction_to_cu_i_20_port, 
                           curr_instruction_to_cu(19) => 
                           curr_instruction_to_cu_i_19_port, 
                           curr_instruction_to_cu(18) => 
                           curr_instruction_to_cu_i_18_port, 
                           curr_instruction_to_cu(17) => 
                           curr_instruction_to_cu_i_17_port, 
                           curr_instruction_to_cu(16) => 
                           curr_instruction_to_cu_i_16_port, 
                           curr_instruction_to_cu(15) => 
                           curr_instruction_to_cu_i_15_port, 
                           curr_instruction_to_cu(14) => 
                           curr_instruction_to_cu_i_14_port, 
                           curr_instruction_to_cu(13) => 
                           curr_instruction_to_cu_i_13_port, 
                           curr_instruction_to_cu(12) => 
                           curr_instruction_to_cu_i_12_port, 
                           curr_instruction_to_cu(11) => 
                           curr_instruction_to_cu_i_11_port, 
                           curr_instruction_to_cu(10) => 
                           curr_instruction_to_cu_i_10_port, 
                           curr_instruction_to_cu(9) => 
                           curr_instruction_to_cu_i_9_port, 
                           curr_instruction_to_cu(8) => 
                           curr_instruction_to_cu_i_8_port, 
                           curr_instruction_to_cu(7) => 
                           curr_instruction_to_cu_i_7_port, 
                           curr_instruction_to_cu(6) => 
                           curr_instruction_to_cu_i_6_port, 
                           curr_instruction_to_cu(5) => 
                           curr_instruction_to_cu_i_5_port, 
                           curr_instruction_to_cu(4) => 
                           curr_instruction_to_cu_i_4_port, 
                           curr_instruction_to_cu(3) => 
                           curr_instruction_to_cu_i_3_port, 
                           curr_instruction_to_cu(2) => 
                           curr_instruction_to_cu_i_2_port, 
                           curr_instruction_to_cu(1) => 
                           curr_instruction_to_cu_i_1_port, 
                           curr_instruction_to_cu(0) => 
                           curr_instruction_to_cu_i_0_port, enable_rf => 
                           enable_rf_i, read_rf_p1 => read_rf_p1_i, read_rf_p2 
                           => read_rf_p2_i, write_rf => write_rf_i, 
                           rtype_itypen => rtype_itypen_i, compute_sext => 
                           compute_sext_i, jump_sext => jump_sext_i, 
                           alu_op_type(3) => alu_op_type_i_3_port, 
                           alu_op_type(2) => alu_op_type_i_2_port, 
                           alu_op_type(1) => alu_op_type_i_1_port, 
                           alu_op_type(0) => alu_op_type_i_0_port, sel_val_a =>
                           sel_val_a_i_0_port, sel_val_b => sel_val_b_i_0_port,
                           signed_notsigned => signed_notsigned_i, 
                           evaluate_branch(1) => evaluate_branch_i_1_port, 
                           evaluate_branch(0) => evaluate_branch_i_0_port, 
                           alu_cin => alu_cin_i, alu_overflow => alu_overflow_i
                           , zero_mul_detect => zero_mul_detect_i, 
                           mul_exeception => mul_exeception_i, dram_enable_cu 
                           => dram_enable_cu_i, dram_r_nw_cu => dram_r_nw_cu_i,
                           dram_ready_cu => dram_ready_cu_i, update_pc_branch 
                           => update_pc_branch_i, select_wb => 
                           select_wb_i_0_port);
   DRAM_ADDRESS_0_port <= '0';

end SYN_dlx_rtl;
